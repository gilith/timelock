/*----------------------------------------------------------------------------+
| module test_timelock_3 satisfies the following property:                    |
|                                                                             |
| !x t.                                                                       |
|     ?d. !j. (!i. i <= d + j ==> (signal ld (t + i) <=> i <= 11)) /\         |
|             (bits_to_num (bsignal xs[0:183] (t + 22)) +                     |
|              2 * bits_to_num (bsignal xc[0:183] (t + 22))) MOD              |
|             (99891253338474858246474952633767320929 * checksum_prime) =     |
|             (x * 2 EXP 186) MOD                                             |
|             (99891253338474858246474952633767320929 * checksum_prime)       |
|             ==> (!i. i <= d + j ==> (signal dn (t + 11 + i) <=> d <= i)) /\ |
|                 (bits_to_num (bsignal ys[0:183] (t + 11 + d + j)) +         |
|                  2 * bits_to_num (bsignal yc[0:183] (t + 11 + d + j))) MOD  |
|                 (99891253338474858246474952633767320929 * checksum_prime) = |
|                 (x EXP (2 EXP (10 EXP 3)) * 2 EXP 186) MOD                  |
|                 (99891253338474858246474952633767320929 * checksum_prime)   |
|                                                                             |
| where checksum_prime = 201301130512090183.                                  |
|                                                                             |
| How to use the module:                                                      |
|                                                                             |
|   1. Hold the ld signal high for at least 12 cycles.                        |
|      Load the input into the xs and xc buses.                               |
|   2. Drop the ld signal low.                                                |
|   3. Wait 208,011 cycles for the dn signal to go high.                      |
|   4. Read the result from the ys and yc buses.                              |
|                                                                             |
| Assuming the circuit is clocked at 1GHz, the above computation will take    |
| ~0.0002 seconds.                                                            |
|                                                                             |
| Copyright (c) 2014 Joe Leslie-Hurd, distributed under the MIT license       |
+----------------------------------------------------------------------------*/

module test_timelock_3(clk,ld,xs,xc,dn,ys,yc);
  input clk;
  input ld;
  input [183:0] xs;
  input [183:0] xc;

  output dn;
  output [183:0] ys;
  output [183:0] yc;

  reg ctre_cp0;  // 3:4|2/1=2
  reg ctre_cp1;  // 4:4|2/1=2
  reg ctre_cp2;  // 4:4|2/1=2
  reg ctre_cp3;  // 4:4|2/1=2
  reg ctre_cp4;  // 4:4|2/1=2
  reg ctre_cp5;  // 4:4|2/1=2
  reg ctre_cp6;  // 4:4|2/1=2
  reg ctre_cp7;  // 4:4|2/1=2
  reg ctre_cp8;  // 4:4|2/1=2
  reg ctre_cp9;  // 4:4|2/1=2
  reg ctre_dp;  // 4:4|2/1=2
  reg ctre_sp0;  // 3:3|2/1=2
  reg ctre_sp1;  // 4:4|2/1=2
  reg ctre_sp2;  // 4:4|2/1=2
  reg ctre_sp3;  // 4:3|2/1=2
  reg ctre_sp4;  // 4:3|2/1=2
  reg ctre_sp5;  // 4:4|2/1=2
  reg ctre_sp6;  // 4:4|2/1=2
  reg ctre_sp7;  // 4:4|2/1=2
  reg ctre_sp8;  // 4:4|2/1=2
  reg ctre_sp9;  // 4:4|2/1=2
  reg multm_compress_ncd;  // 1:0|248/54=4
  reg multm_compress_nsd;  // 1:0|278/60=4
  reg multm_compress_pipe0_x1;  // 2:1|1/1=1
  reg multm_compress_pipe0_x2;  // 1:0|1/1=3
  reg multm_compress_pipe0_x3;  // 1:0|1/3=4
  reg multm_compress_pipe0_x4;  // 1:0|1/13=4
  reg multm_compress_pipe1_x1;  // 3:2|1/1=1
  reg multm_compress_pipe1_x2;  // 1:0|1/1=3
  reg multm_compress_pipe1_x3;  // 1:0|1/3=4
  reg multm_compress_pipe1_x4;  // 1:0|1/12=4
  reg multm_ctrp_ctr_cp0;  // 2:2|3/1=3
  reg multm_ctrp_ctr_cp1;  // 3:3|2/1=2
  reg multm_ctrp_ctr_cp2;  // 3:3|2/1=2
  reg multm_ctrp_ctr_cp3;  // 3:3|2/1=2
  reg multm_ctrp_ctr_cp4;  // 3:3|2/1=2
  reg multm_ctrp_ctr_cp5;  // 3:3|2/1=2
  reg multm_ctrp_ctr_cp6;  // 3:3|2/1=2
  reg multm_ctrp_ctr_cp7;  // 3:3|4/1=4
  reg multm_ctrp_ctr_dp;  // 3:3|4/1=4
  reg multm_ctrp_ctr_sp0;  // 3:2|2/1=2
  reg multm_ctrp_ctr_sp1;  // 3:3|2/1=2
  reg multm_ctrp_ctr_sp2;  // 3:3|2/1=2
  reg multm_ctrp_ctr_sp3;  // 3:3|2/1=2
  reg multm_ctrp_ctr_sp4;  // 3:3|2/1=2
  reg multm_ctrp_ctr_sp5;  // 3:2|2/1=2
  reg multm_ctrp_ctr_sp6;  // 3:3|2/1=2
  reg multm_jpd;  // 1:0|370/71=5
  reg multm_pipe_x1;  // 3:5|1/1=1
  reg multm_pipe_x2;  // 1:0|1/1=3
  reg multm_pipe_x3;  // 1:0|1/3=4
  reg multm_pipe_x4;  // 1:0|1/14=5
  reg multm_qcp0;  // 5:6|3/1=3
  reg multm_qcp1;  // 5:6|3/1=3
  reg multm_qcp2;  // 5:6|3/1=3
  reg multm_qcp3;  // 5:6|3/1=3
  reg multm_qcp4;  // 5:6|3/1=3
  reg multm_qcp5;  // 5:6|3/1=3
  reg multm_qcp6;  // 5:6|3/1=3
  reg multm_qcp7;  // 5:6|3/1=3
  reg multm_qcp8;  // 5:6|3/1=3
  reg multm_qcp9;  // 5:6|3/1=3
  reg multm_qcp10;  // 2:2|3/1=3
  reg multm_qcp11;  // 9:13|3/1=3
  reg multm_qcp12;  // 9:13|3/1=3
  reg multm_qcp13;  // 9:13|3/1=3
  reg multm_qcp14;  // 9:13|3/1=3
  reg multm_qcp15;  // 9:13|3/1=3
  reg multm_qcp16;  // 9:13|3/1=3
  reg multm_qcp17;  // 9:13|3/1=3
  reg multm_qcp18;  // 9:13|3/1=3
  reg multm_qcp19;  // 9:13|3/1=3
  reg multm_qcp20;  // 9:13|3/1=3
  reg multm_qcp21;  // 9:13|3/1=3
  reg multm_qcp22;  // 9:13|3/1=3
  reg multm_qcp23;  // 9:13|3/1=3
  reg multm_qcp24;  // 9:13|3/1=3
  reg multm_qcp25;  // 9:13|3/1=3
  reg multm_qcp26;  // 9:13|3/1=3
  reg multm_qcp27;  // 9:13|3/1=3
  reg multm_qcp28;  // 9:13|3/1=3
  reg multm_qcp29;  // 9:13|3/1=3
  reg multm_qcp30;  // 9:13|3/1=3
  reg multm_qcp31;  // 9:13|3/1=3
  reg multm_qcp32;  // 9:13|3/1=3
  reg multm_qcp33;  // 9:13|3/1=3
  reg multm_qcp34;  // 9:13|3/1=3
  reg multm_qcp35;  // 9:13|3/1=3
  reg multm_qcp36;  // 9:13|3/1=3
  reg multm_qcp37;  // 9:13|3/1=3
  reg multm_qcp38;  // 9:13|3/1=3
  reg multm_qcp39;  // 9:13|3/1=3
  reg multm_qcp40;  // 9:13|3/1=3
  reg multm_qcp41;  // 9:13|3/1=3
  reg multm_qcp42;  // 9:13|3/1=3
  reg multm_qcp43;  // 9:13|3/1=3
  reg multm_qcp44;  // 9:13|3/1=3
  reg multm_qcp45;  // 9:13|3/1=3
  reg multm_qcp46;  // 9:13|3/1=3
  reg multm_qcp47;  // 9:13|3/1=3
  reg multm_qcp48;  // 9:13|3/1=3
  reg multm_qcp49;  // 9:13|3/1=3
  reg multm_qcp50;  // 9:13|3/1=3
  reg multm_qcp51;  // 9:13|3/1=3
  reg multm_qcp52;  // 9:13|3/1=3
  reg multm_qcp53;  // 9:13|3/1=3
  reg multm_qcp54;  // 9:13|3/1=3
  reg multm_qcp55;  // 9:13|3/1=3
  reg multm_qcp56;  // 9:13|3/1=3
  reg multm_qcp57;  // 9:13|3/1=3
  reg multm_qcp58;  // 9:13|3/1=3
  reg multm_qcp59;  // 9:13|3/1=3
  reg multm_qcp60;  // 9:13|3/1=3
  reg multm_qcp61;  // 9:13|3/1=3
  reg multm_qcp62;  // 9:13|3/1=3
  reg multm_qcp63;  // 9:13|3/1=3
  reg multm_qcp64;  // 9:13|3/1=3
  reg multm_qcp65;  // 9:13|3/1=3
  reg multm_qcp66;  // 9:13|3/1=3
  reg multm_qcp67;  // 9:13|3/1=3
  reg multm_qcp68;  // 9:13|3/1=3
  reg multm_qcp69;  // 9:13|3/1=3
  reg multm_qcp70;  // 9:13|3/1=3
  reg multm_qcp71;  // 9:13|3/1=3
  reg multm_qcp72;  // 9:13|3/1=3
  reg multm_qcp73;  // 9:13|3/1=3
  reg multm_qcp74;  // 9:13|3/1=3
  reg multm_qcp75;  // 9:13|3/1=3
  reg multm_qcp76;  // 9:13|3/1=3
  reg multm_qcp77;  // 9:13|3/1=3
  reg multm_qcp78;  // 9:13|3/1=3
  reg multm_qcp79;  // 9:13|3/1=3
  reg multm_qcp80;  // 9:13|3/1=3
  reg multm_qcp81;  // 9:13|3/1=3
  reg multm_qcp82;  // 9:13|3/1=3
  reg multm_qcp83;  // 9:13|3/1=3
  reg multm_qcp84;  // 9:13|3/1=3
  reg multm_qcp85;  // 9:13|3/1=3
  reg multm_qcp86;  // 9:13|3/1=3
  reg multm_qcp87;  // 9:13|3/1=3
  reg multm_qcp88;  // 9:13|3/1=3
  reg multm_qcp89;  // 9:13|3/1=3
  reg multm_qcp90;  // 9:13|3/1=3
  reg multm_qcp91;  // 9:13|3/1=3
  reg multm_qcp92;  // 9:13|3/1=3
  reg multm_qcp93;  // 9:13|3/1=3
  reg multm_qcp94;  // 9:13|3/1=3
  reg multm_qcp95;  // 9:13|3/1=3
  reg multm_qcp96;  // 9:13|3/1=3
  reg multm_qcp97;  // 9:13|3/1=3
  reg multm_qcp98;  // 9:13|3/1=3
  reg multm_qcp99;  // 9:13|3/1=3
  reg multm_qcp100;  // 9:13|3/1=3
  reg multm_qcp101;  // 9:13|3/1=3
  reg multm_qcp102;  // 9:13|3/1=3
  reg multm_qcp103;  // 9:13|3/1=3
  reg multm_qcp104;  // 9:13|3/1=3
  reg multm_qcp105;  // 9:13|3/1=3
  reg multm_qcp106;  // 9:13|3/1=3
  reg multm_qcp107;  // 9:13|3/1=3
  reg multm_qcp108;  // 9:13|3/1=3
  reg multm_qcp109;  // 9:13|3/1=3
  reg multm_qcp110;  // 9:13|3/1=3
  reg multm_qcp111;  // 9:13|3/1=3
  reg multm_qcp112;  // 9:13|3/1=3
  reg multm_qcp113;  // 9:13|3/1=3
  reg multm_qcp114;  // 9:13|3/1=3
  reg multm_qcp115;  // 9:13|3/1=3
  reg multm_qcp116;  // 9:13|3/1=3
  reg multm_qcp117;  // 9:13|3/1=3
  reg multm_qcp118;  // 9:13|3/1=3
  reg multm_qcp119;  // 9:13|3/1=3
  reg multm_qcp120;  // 9:13|3/1=3
  reg multm_qcp121;  // 9:13|3/1=3
  reg multm_qcp122;  // 9:13|3/1=3
  reg multm_qcp123;  // 9:13|3/1=3
  reg multm_qcp124;  // 9:13|3/1=3
  reg multm_qcp125;  // 9:13|3/1=3
  reg multm_qcp126;  // 9:13|3/1=3
  reg multm_qcp127;  // 9:13|3/1=3
  reg multm_qcp128;  // 9:13|3/1=3
  reg multm_qcp129;  // 9:13|3/1=3
  reg multm_qcp130;  // 9:13|3/1=3
  reg multm_qcp131;  // 9:13|3/1=3
  reg multm_qcp132;  // 9:13|3/1=3
  reg multm_qcp133;  // 9:13|3/1=3
  reg multm_qcp134;  // 9:13|3/1=3
  reg multm_qcp135;  // 9:13|3/1=3
  reg multm_qcp136;  // 9:13|3/1=3
  reg multm_qcp137;  // 9:13|3/1=3
  reg multm_qcp138;  // 9:13|3/1=3
  reg multm_qcp139;  // 9:13|3/1=3
  reg multm_qcp140;  // 9:13|3/1=3
  reg multm_qcp141;  // 9:13|3/1=3
  reg multm_qcp142;  // 9:13|3/1=3
  reg multm_qcp143;  // 9:13|3/1=3
  reg multm_qcp144;  // 9:13|3/1=3
  reg multm_qcp145;  // 9:13|3/1=3
  reg multm_qcp146;  // 9:13|3/1=3
  reg multm_qcp147;  // 9:13|3/1=3
  reg multm_qcp148;  // 9:13|3/1=3
  reg multm_qcp149;  // 9:13|3/1=3
  reg multm_qcp150;  // 9:13|3/1=3
  reg multm_qcp151;  // 9:13|3/1=3
  reg multm_qcp152;  // 9:13|3/1=3
  reg multm_qcp153;  // 9:13|3/1=3
  reg multm_qcp154;  // 9:13|3/1=3
  reg multm_qcp155;  // 9:13|3/1=3
  reg multm_qcp156;  // 9:13|3/1=3
  reg multm_qcp157;  // 9:13|3/1=3
  reg multm_qcp158;  // 9:13|3/1=3
  reg multm_qcp159;  // 9:13|3/1=3
  reg multm_qcp160;  // 9:13|3/1=3
  reg multm_qcp161;  // 9:13|3/1=3
  reg multm_qcp162;  // 9:13|3/1=3
  reg multm_qcp163;  // 9:13|3/1=3
  reg multm_qcp164;  // 9:13|3/1=3
  reg multm_qcp165;  // 9:13|3/1=3
  reg multm_qcp166;  // 9:13|3/1=3
  reg multm_qcp167;  // 9:13|3/1=3
  reg multm_qcp168;  // 9:13|3/1=3
  reg multm_qcp169;  // 9:13|3/1=3
  reg multm_qcp170;  // 9:13|3/1=3
  reg multm_qcp171;  // 9:13|3/1=3
  reg multm_qcp172;  // 9:13|3/1=3
  reg multm_qcp173;  // 9:13|3/1=3
  reg multm_qcp174;  // 9:13|3/1=3
  reg multm_qcp175;  // 9:13|3/1=3
  reg multm_qcp176;  // 9:13|3/1=3
  reg multm_qcp177;  // 9:13|3/1=3
  reg multm_qcp178;  // 9:13|3/1=3
  reg multm_qcp179;  // 9:13|3/1=3
  reg multm_qcp180;  // 9:13|3/1=3
  reg multm_qcp181;  // 9:13|3/1=3
  reg multm_qcp182;  // 9:13|3/1=3
  reg multm_qcp183;  // 8:12|3/1=3
  reg multm_qcp184;  // 8:9|2/1=2
  reg multm_qsp0;  // 5:3|3/1=3
  reg multm_qsp1;  // 5:3|3/1=3
  reg multm_qsp2;  // 5:3|3/1=3
  reg multm_qsp3;  // 5:3|3/1=3
  reg multm_qsp4;  // 5:3|3/1=3
  reg multm_qsp5;  // 5:3|3/1=3
  reg multm_qsp6;  // 5:3|3/1=3
  reg multm_qsp7;  // 5:3|3/1=3
  reg multm_qsp8;  // 5:3|3/1=3
  reg multm_qsp9;  // 5:3|3/1=3
  reg multm_qsp10;  // 5:3|3/1=3
  reg multm_qsp11;  // 9:10|3/1=3
  reg multm_qsp12;  // 9:10|3/1=3
  reg multm_qsp13;  // 9:10|3/1=3
  reg multm_qsp14;  // 9:10|3/1=3
  reg multm_qsp15;  // 9:10|3/1=3
  reg multm_qsp16;  // 9:10|3/1=3
  reg multm_qsp17;  // 9:10|3/1=3
  reg multm_qsp18;  // 9:10|3/1=3
  reg multm_qsp19;  // 9:10|3/1=3
  reg multm_qsp20;  // 9:10|3/1=3
  reg multm_qsp21;  // 9:10|3/1=3
  reg multm_qsp22;  // 9:10|3/1=3
  reg multm_qsp23;  // 9:10|3/1=3
  reg multm_qsp24;  // 9:10|3/1=3
  reg multm_qsp25;  // 9:10|3/1=3
  reg multm_qsp26;  // 9:10|3/1=3
  reg multm_qsp27;  // 9:10|3/1=3
  reg multm_qsp28;  // 9:10|3/1=3
  reg multm_qsp29;  // 9:10|3/1=3
  reg multm_qsp30;  // 9:10|3/1=3
  reg multm_qsp31;  // 9:10|3/1=3
  reg multm_qsp32;  // 9:10|3/1=3
  reg multm_qsp33;  // 9:10|3/1=3
  reg multm_qsp34;  // 9:10|3/1=3
  reg multm_qsp35;  // 9:10|3/1=3
  reg multm_qsp36;  // 9:10|3/1=3
  reg multm_qsp37;  // 9:10|3/1=3
  reg multm_qsp38;  // 9:10|3/1=3
  reg multm_qsp39;  // 9:10|3/1=3
  reg multm_qsp40;  // 9:10|3/1=3
  reg multm_qsp41;  // 9:10|3/1=3
  reg multm_qsp42;  // 9:10|3/1=3
  reg multm_qsp43;  // 9:10|3/1=3
  reg multm_qsp44;  // 9:10|3/1=3
  reg multm_qsp45;  // 9:10|3/1=3
  reg multm_qsp46;  // 9:10|3/1=3
  reg multm_qsp47;  // 9:10|3/1=3
  reg multm_qsp48;  // 9:10|3/1=3
  reg multm_qsp49;  // 9:10|3/1=3
  reg multm_qsp50;  // 9:10|3/1=3
  reg multm_qsp51;  // 9:10|3/1=3
  reg multm_qsp52;  // 9:10|3/1=3
  reg multm_qsp53;  // 9:10|3/1=3
  reg multm_qsp54;  // 9:10|3/1=3
  reg multm_qsp55;  // 9:10|3/1=3
  reg multm_qsp56;  // 9:10|3/1=3
  reg multm_qsp57;  // 9:10|3/1=3
  reg multm_qsp58;  // 9:10|3/1=3
  reg multm_qsp59;  // 9:10|3/1=3
  reg multm_qsp60;  // 9:10|3/1=3
  reg multm_qsp61;  // 9:10|3/1=3
  reg multm_qsp62;  // 9:10|3/1=3
  reg multm_qsp63;  // 9:10|3/1=3
  reg multm_qsp64;  // 9:10|3/1=3
  reg multm_qsp65;  // 9:10|3/1=3
  reg multm_qsp66;  // 9:10|3/1=3
  reg multm_qsp67;  // 9:10|3/1=3
  reg multm_qsp68;  // 9:10|3/1=3
  reg multm_qsp69;  // 9:10|3/1=3
  reg multm_qsp70;  // 9:10|3/1=3
  reg multm_qsp71;  // 9:10|3/1=3
  reg multm_qsp72;  // 9:10|3/1=3
  reg multm_qsp73;  // 9:10|3/1=3
  reg multm_qsp74;  // 9:10|3/1=3
  reg multm_qsp75;  // 9:10|3/1=3
  reg multm_qsp76;  // 9:10|3/1=3
  reg multm_qsp77;  // 9:10|3/1=3
  reg multm_qsp78;  // 9:10|3/1=3
  reg multm_qsp79;  // 9:10|3/1=3
  reg multm_qsp80;  // 9:10|3/1=3
  reg multm_qsp81;  // 9:10|3/1=3
  reg multm_qsp82;  // 9:10|3/1=3
  reg multm_qsp83;  // 9:10|3/1=3
  reg multm_qsp84;  // 9:10|3/1=3
  reg multm_qsp85;  // 9:10|3/1=3
  reg multm_qsp86;  // 9:10|3/1=3
  reg multm_qsp87;  // 9:10|3/1=3
  reg multm_qsp88;  // 9:10|3/1=3
  reg multm_qsp89;  // 9:10|3/1=3
  reg multm_qsp90;  // 9:10|3/1=3
  reg multm_qsp91;  // 9:10|3/1=3
  reg multm_qsp92;  // 9:10|3/1=3
  reg multm_qsp93;  // 9:10|3/1=3
  reg multm_qsp94;  // 9:10|3/1=3
  reg multm_qsp95;  // 9:10|3/1=3
  reg multm_qsp96;  // 9:10|3/1=3
  reg multm_qsp97;  // 9:10|3/1=3
  reg multm_qsp98;  // 9:10|3/1=3
  reg multm_qsp99;  // 9:10|3/1=3
  reg multm_qsp100;  // 9:10|3/1=3
  reg multm_qsp101;  // 9:10|3/1=3
  reg multm_qsp102;  // 9:10|3/1=3
  reg multm_qsp103;  // 9:10|3/1=3
  reg multm_qsp104;  // 9:10|3/1=3
  reg multm_qsp105;  // 9:10|3/1=3
  reg multm_qsp106;  // 9:10|3/1=3
  reg multm_qsp107;  // 9:10|3/1=3
  reg multm_qsp108;  // 9:10|3/1=3
  reg multm_qsp109;  // 9:10|3/1=3
  reg multm_qsp110;  // 9:10|3/1=3
  reg multm_qsp111;  // 9:10|3/1=3
  reg multm_qsp112;  // 9:10|3/1=3
  reg multm_qsp113;  // 9:10|3/1=3
  reg multm_qsp114;  // 9:10|3/1=3
  reg multm_qsp115;  // 9:10|3/1=3
  reg multm_qsp116;  // 9:10|3/1=3
  reg multm_qsp117;  // 9:10|3/1=3
  reg multm_qsp118;  // 9:10|3/1=3
  reg multm_qsp119;  // 9:10|3/1=3
  reg multm_qsp120;  // 9:10|3/1=3
  reg multm_qsp121;  // 9:10|3/1=3
  reg multm_qsp122;  // 9:10|3/1=3
  reg multm_qsp123;  // 9:10|3/1=3
  reg multm_qsp124;  // 9:10|3/1=3
  reg multm_qsp125;  // 9:10|3/1=3
  reg multm_qsp126;  // 9:10|3/1=3
  reg multm_qsp127;  // 9:10|3/1=3
  reg multm_qsp128;  // 9:10|3/1=3
  reg multm_qsp129;  // 9:10|3/1=3
  reg multm_qsp130;  // 9:10|3/1=3
  reg multm_qsp131;  // 9:10|3/1=3
  reg multm_qsp132;  // 9:10|3/1=3
  reg multm_qsp133;  // 9:10|3/1=3
  reg multm_qsp134;  // 9:10|3/1=3
  reg multm_qsp135;  // 9:10|3/1=3
  reg multm_qsp136;  // 9:10|3/1=3
  reg multm_qsp137;  // 9:10|3/1=3
  reg multm_qsp138;  // 9:10|3/1=3
  reg multm_qsp139;  // 9:10|3/1=3
  reg multm_qsp140;  // 9:10|3/1=3
  reg multm_qsp141;  // 9:10|3/1=3
  reg multm_qsp142;  // 9:10|3/1=3
  reg multm_qsp143;  // 9:10|3/1=3
  reg multm_qsp144;  // 9:10|3/1=3
  reg multm_qsp145;  // 9:10|3/1=3
  reg multm_qsp146;  // 9:10|3/1=3
  reg multm_qsp147;  // 9:10|3/1=3
  reg multm_qsp148;  // 9:10|3/1=3
  reg multm_qsp149;  // 9:10|3/1=3
  reg multm_qsp150;  // 9:10|3/1=3
  reg multm_qsp151;  // 9:10|3/1=3
  reg multm_qsp152;  // 9:10|3/1=3
  reg multm_qsp153;  // 9:10|3/1=3
  reg multm_qsp154;  // 9:10|3/1=3
  reg multm_qsp155;  // 9:10|3/1=3
  reg multm_qsp156;  // 9:10|3/1=3
  reg multm_qsp157;  // 9:10|3/1=3
  reg multm_qsp158;  // 9:10|3/1=3
  reg multm_qsp159;  // 9:10|3/1=3
  reg multm_qsp160;  // 9:10|3/1=3
  reg multm_qsp161;  // 9:10|3/1=3
  reg multm_qsp162;  // 9:10|3/1=3
  reg multm_qsp163;  // 9:10|3/1=3
  reg multm_qsp164;  // 9:10|3/1=3
  reg multm_qsp165;  // 9:10|3/1=3
  reg multm_qsp166;  // 9:10|3/1=3
  reg multm_qsp167;  // 9:10|3/1=3
  reg multm_qsp168;  // 9:10|3/1=3
  reg multm_qsp169;  // 9:10|3/1=3
  reg multm_qsp170;  // 9:10|3/1=3
  reg multm_qsp171;  // 9:10|3/1=3
  reg multm_qsp172;  // 9:10|3/1=3
  reg multm_qsp173;  // 9:10|3/1=3
  reg multm_qsp174;  // 9:10|3/1=3
  reg multm_qsp175;  // 9:10|3/1=3
  reg multm_qsp176;  // 9:10|3/1=3
  reg multm_qsp177;  // 9:10|3/1=3
  reg multm_qsp178;  // 9:10|3/1=3
  reg multm_qsp179;  // 9:10|3/1=3
  reg multm_qsp180;  // 9:10|3/1=3
  reg multm_qsp181;  // 9:10|3/1=3
  reg multm_qsp182;  // 9:10|3/1=3
  reg multm_qsp183;  // 8:9|3/1=3
  reg multm_qsp184;  // 6:4|3/1=3
  reg multm_reduce_ld1;  // 1:0|372/72=5
  reg multm_reduce_ld2;  // 1:0|367/71=5
  reg multm_reduce_mulb0_cp0;  // 5:7|4/1=4
  reg multm_reduce_mulb0_cp1;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp2;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp3;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp4;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp5;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp6;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp7;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp8;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp9;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp10;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp11;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp12;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp13;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp14;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp15;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp16;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp17;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp18;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp19;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp20;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp21;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp22;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp23;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp24;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp25;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp26;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp27;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp28;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp29;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp30;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp31;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp32;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp33;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp34;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp35;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp36;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp37;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp38;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp39;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp40;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp41;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp42;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp43;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp44;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp45;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp46;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp47;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp48;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp49;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp50;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp51;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp52;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp53;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp54;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp55;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp56;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp57;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp58;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp59;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp60;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp61;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp62;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp63;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp64;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp65;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp66;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp67;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp68;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp69;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp70;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp71;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp72;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp73;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp74;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp75;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp76;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp77;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp78;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp79;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp80;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp81;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp82;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp83;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp84;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp85;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp86;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp87;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp88;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp89;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp90;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp91;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp92;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp93;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp94;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp95;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp96;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp97;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp98;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp99;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp100;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp101;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp102;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp103;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp104;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp105;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp106;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp107;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp108;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp109;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp110;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp111;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp112;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp113;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp114;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp115;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp116;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp117;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp118;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp119;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp120;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp121;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp122;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp123;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp124;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp125;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp126;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp127;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp128;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp129;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp130;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp131;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp132;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp133;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp134;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp135;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp136;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp137;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp138;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp139;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp140;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp141;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp142;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp143;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp144;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp145;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp146;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp147;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp148;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp149;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp150;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp151;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp152;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp153;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp154;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp155;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp156;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp157;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp158;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp159;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp160;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp161;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp162;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp163;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp164;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp165;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp166;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp167;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp168;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp169;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp170;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp171;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp172;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp173;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp174;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp175;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp176;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp177;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp178;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp179;  // 6:12|4/1=4
  reg multm_reduce_mulb0_cp180;  // 5:8|4/1=4
  reg multm_reduce_mulb0_cp181;  // 6:9|4/1=4
  reg multm_reduce_mulb0_cp182;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp183;  // 6:13|4/1=4
  reg multm_reduce_mulb0_cp184;  // 5:14|2/1=2
  reg multm_reduce_mulb0_sp0;  // 5:7|3/1=3
  reg multm_reduce_mulb0_sp1;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp2;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp3;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp4;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp5;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp6;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp7;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp8;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp9;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp10;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp11;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp12;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp13;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp14;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp15;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp16;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp17;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp18;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp19;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp20;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp21;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp22;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp23;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp24;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp25;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp26;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp27;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp28;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp29;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp30;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp31;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp32;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp33;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp34;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp35;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp36;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp37;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp38;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp39;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp40;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp41;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp42;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp43;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp44;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp45;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp46;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp47;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp48;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp49;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp50;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp51;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp52;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp53;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp54;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp55;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp56;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp57;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp58;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp59;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp60;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp61;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp62;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp63;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp64;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp65;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp66;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp67;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp68;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp69;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp70;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp71;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp72;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp73;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp74;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp75;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp76;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp77;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp78;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp79;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp80;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp81;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp82;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp83;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp84;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp85;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp86;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp87;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp88;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp89;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp90;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp91;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp92;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp93;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp94;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp95;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp96;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp97;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp98;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp99;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp100;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp101;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp102;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp103;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp104;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp105;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp106;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp107;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp108;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp109;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp110;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp111;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp112;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp113;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp114;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp115;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp116;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp117;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp118;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp119;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp120;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp121;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp122;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp123;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp124;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp125;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp126;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp127;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp128;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp129;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp130;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp131;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp132;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp133;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp134;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp135;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp136;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp137;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp138;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp139;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp140;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp141;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp142;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp143;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp144;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp145;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp146;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp147;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp148;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp149;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp150;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp151;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp152;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp153;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp154;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp155;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp156;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp157;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp158;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp159;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp160;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp161;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp162;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp163;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp164;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp165;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp166;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp167;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp168;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp169;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp170;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp171;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp172;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp173;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp174;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp175;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp176;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp177;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp178;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp179;  // 6:12|4/1=4
  reg multm_reduce_mulb0_sp180;  // 5:8|4/1=4
  reg multm_reduce_mulb0_sp181;  // 6:9|4/1=4
  reg multm_reduce_mulb0_sp182;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp183;  // 6:13|4/1=4
  reg multm_reduce_mulb0_sp184;  // 5:11|4/1=4
  reg multm_reduce_mulsc_mulb_cp175;  // 9:20|4/1=4
  reg multm_reduce_mulsc_mulb_cp176;  // 9:20|4/1=4
  reg multm_reduce_mulsc_mulb_cp177;  // 9:20|4/1=4
  reg multm_reduce_mulsc_mulb_cp178;  // 9:20|4/1=4
  reg multm_reduce_mulsc_mulb_cp179;  // 9:20|4/1=4
  reg multm_reduce_mulsc_mulb_cp180;  // 9:20|4/1=4
  reg multm_reduce_mulsc_mulb_cp181;  // 9:20|4/1=4
  reg multm_reduce_mulsc_mulb_cp182;  // 9:20|4/1=4
  reg multm_reduce_mulsc_mulb_cp183;  // 7:16|2/1=2
  reg multm_reduce_mulsc_mulb_sp176;  // 9:17|4/1=4
  reg multm_reduce_mulsc_mulb_sp177;  // 9:17|4/1=4
  reg multm_reduce_mulsc_mulb_sp178;  // 9:17|4/1=4
  reg multm_reduce_mulsc_mulb_sp179;  // 9:17|4/1=4
  reg multm_reduce_mulsc_mulb_sp180;  // 9:17|4/1=4
  reg multm_reduce_mulsc_mulb_sp181;  // 9:17|4/1=4
  reg multm_reduce_mulsc_mulb_sp182;  // 9:17|4/1=4
  reg multm_reduce_mulsc_mulb_sp183;  // 7:13|4/1=4
  reg multm_reduce_mulsc_pipe_x1;  // 4:2|1/1=1
  reg multm_reduce_mulsc_pipe_x2;  // 1:0|1/1=3
  reg multm_reduce_mulsc_pipe_x3;  // 1:0|1/3=4
  reg multm_reduce_mulsc_pipe_x4;  // 1:0|1/14=5
  reg multm_reduce_mulsc_shrsc_cp0;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp1;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp2;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp3;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp4;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp5;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp6;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp7;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp8;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp9;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp10;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp11;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp12;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp13;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp14;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp15;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp16;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp17;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp18;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp19;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp20;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp21;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp22;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp23;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp24;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp25;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp26;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp27;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp28;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp29;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp30;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp31;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp32;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp33;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp34;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp35;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp36;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp37;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp38;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp39;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp40;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp41;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp42;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp43;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp44;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp45;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp46;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp47;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp48;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp49;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp50;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp51;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp52;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp53;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp54;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp55;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp56;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp57;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp58;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp59;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp60;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp61;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp62;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp63;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp64;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp65;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp66;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp67;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp68;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp69;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp70;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp71;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp72;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp73;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp74;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp75;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp76;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp77;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp78;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp79;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp80;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp81;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp82;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp83;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp84;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp85;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp86;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp87;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp88;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp89;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp90;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp91;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp92;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp93;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp94;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp95;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp96;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp97;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp98;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp99;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp100;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp101;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp102;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp103;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp104;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp105;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp106;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp107;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp108;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp109;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp110;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp111;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp112;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp113;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp114;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp115;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp116;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp117;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp118;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp119;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp120;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp121;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp122;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp123;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp124;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp125;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp126;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp127;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp128;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp129;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp130;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp131;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp132;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp133;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp134;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp135;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp136;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp137;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp138;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp139;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp140;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp141;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp142;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp143;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp144;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp145;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp146;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp147;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp148;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp149;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp150;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp151;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp152;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp153;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp154;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp155;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp156;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp157;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp158;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp159;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp160;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp161;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp162;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp163;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp164;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp165;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp166;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp167;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp168;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp169;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp170;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp171;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp172;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp173;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp174;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp175;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp176;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp177;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp178;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp179;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp180;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp181;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp182;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_cp183;  // 2:1|1/1=1
  reg multm_reduce_mulsc_shrsc_sp0;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp1;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp2;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp3;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp4;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp5;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp6;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp7;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp8;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp9;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp10;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp11;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp12;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp13;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp14;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp15;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp16;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp17;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp18;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp19;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp20;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp21;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp22;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp23;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp24;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp25;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp26;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp27;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp28;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp29;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp30;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp31;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp32;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp33;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp34;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp35;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp36;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp37;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp38;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp39;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp40;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp41;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp42;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp43;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp44;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp45;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp46;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp47;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp48;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp49;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp50;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp51;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp52;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp53;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp54;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp55;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp56;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp57;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp58;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp59;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp60;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp61;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp62;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp63;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp64;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp65;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp66;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp67;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp68;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp69;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp70;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp71;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp72;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp73;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp74;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp75;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp76;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp77;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp78;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp79;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp80;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp81;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp82;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp83;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp84;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp85;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp86;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp87;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp88;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp89;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp90;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp91;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp92;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp93;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp94;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp95;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp96;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp97;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp98;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp99;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp100;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp101;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp102;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp103;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp104;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp105;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp106;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp107;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp108;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp109;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp110;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp111;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp112;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp113;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp114;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp115;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp116;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp117;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp118;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp119;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp120;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp121;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp122;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp123;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp124;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp125;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp126;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp127;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp128;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp129;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp130;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp131;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp132;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp133;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp134;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp135;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp136;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp137;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp138;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp139;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp140;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp141;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp142;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp143;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp144;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp145;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp146;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp147;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp148;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp149;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp150;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp151;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp152;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp153;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp154;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp155;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp156;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp157;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp158;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp159;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp160;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp161;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp162;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp163;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp164;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp165;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp166;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp167;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp168;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp169;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp170;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp171;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp172;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp173;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp174;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp175;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp176;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp177;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp178;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp179;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp180;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp181;  // 4:2|2/1=2
  reg multm_reduce_mulsc_shrsc_sp182;  // 3:1|2/1=2
  reg multm_reduce_mulsc_xbd;  // 1:0|369/71=5
  reg multm_reduce_pipe0_x1;  // 1:0|1/1=1
  reg multm_reduce_pipe0_x2;  // 1:0|1/1=3
  reg multm_reduce_pipe0_x3;  // 1:0|1/3=4
  reg multm_reduce_pipe0_x4;  // 1:0|1/14=5
  reg multm_reduce_pipe0_x5;  // 1:0|370/71=5
  reg multm_reduce_pipe0_x6;  // 1:0|1/1=1
  reg multm_reduce_pipe0_x7;  // 1:0|1/1=3
  reg multm_reduce_pipe0_x8;  // 1:0|1/3=4
  reg multm_reduce_pipe0_x9;  // 1:0|1/14=5
  reg multm_reduce_pipe1_x1;  // 1:0|1/1=1
  reg multm_reduce_pipe1_x2;  // 1:0|1/1=3
  reg multm_reduce_pipe1_x3;  // 1:0|1/3=4
  reg multm_reduce_pipe1_x4;  // 1:0|1/14=5
  reg multm_reduce_pipe2_x1;  // 3:3|1/1=1
  reg multm_reduce_pipe2_x2;  // 1:0|1/1=3
  reg multm_reduce_pipe2_x3;  // 1:0|1/3=4
  reg multm_reduce_pipe2_x4;  // 1:0|1/13=4
  reg multm_reduce_qb2;  // 1:0|281/60=4
  reg multm_reduce_sa0;  // 1:0|2/1=2
  reg multm_reduce_sa1;  // 1:0|3/1=3
  reg multm_reduce_sa2;  // 1:0|3/1=3
  reg multm_reduce_sa3;  // 1:0|3/1=3
  reg multm_reduce_sa4;  // 1:0|3/1=3
  reg multm_reduce_sa5;  // 1:0|290/37=7
  reg multm_reduce_sa6;  // 1:0|3/5=7
  reg multm_reduce_sa7;  // 1:0|3/1=7
  reg multm_reduce_sa8;  // 1:0|3/1=3
  reg multm_reduce_sa9;  // 4:4|3/1=3
  reg multm_reduce_sa10;  // 8:12|6/1=6
  reg multm_reduce_sa11;  // 9:17|8/1=8
  reg multm_reduce_sa12;  // 9:17|8/1=8
  reg multm_reduce_sa13;  // 9:17|8/1=8
  reg multm_reduce_sa14;  // 9:17|8/1=8
  reg multm_reduce_sa15;  // 9:17|8/1=8
  reg multm_reduce_sa16;  // 9:17|8/1=8
  reg multm_reduce_sa17;  // 9:17|8/1=8
  reg multm_reduce_sa18;  // 9:17|8/1=8
  reg multm_reduce_sa19;  // 9:17|8/1=8
  reg multm_reduce_sa20;  // 9:17|8/1=8
  reg multm_reduce_sa21;  // 9:17|8/1=8
  reg multm_reduce_sa22;  // 9:17|8/1=8
  reg multm_reduce_sa23;  // 9:17|8/1=8
  reg multm_reduce_sa24;  // 9:17|8/1=8
  reg multm_reduce_sa25;  // 9:17|8/1=8
  reg multm_reduce_sa26;  // 9:17|8/1=8
  reg multm_reduce_sa27;  // 9:17|8/1=8
  reg multm_reduce_sa28;  // 9:17|8/1=8
  reg multm_reduce_sa29;  // 9:17|8/1=8
  reg multm_reduce_sa30;  // 9:17|8/1=8
  reg multm_reduce_sa31;  // 9:17|8/1=8
  reg multm_reduce_sa32;  // 9:17|8/1=8
  reg multm_reduce_sa33;  // 9:17|8/1=8
  reg multm_reduce_sa34;  // 9:17|8/1=8
  reg multm_reduce_sa35;  // 9:17|8/1=8
  reg multm_reduce_sa36;  // 9:17|8/1=8
  reg multm_reduce_sa37;  // 9:17|8/1=8
  reg multm_reduce_sa38;  // 9:17|8/1=8
  reg multm_reduce_sa39;  // 9:17|8/1=8
  reg multm_reduce_sa40;  // 9:17|8/1=8
  reg multm_reduce_sa41;  // 9:17|8/1=8
  reg multm_reduce_sa42;  // 9:17|8/1=8
  reg multm_reduce_sa43;  // 9:17|8/1=8
  reg multm_reduce_sa44;  // 9:17|8/1=8
  reg multm_reduce_sa45;  // 9:17|8/1=8
  reg multm_reduce_sa46;  // 9:17|8/1=8
  reg multm_reduce_sa47;  // 9:17|8/1=8
  reg multm_reduce_sa48;  // 9:17|8/1=8
  reg multm_reduce_sa49;  // 9:17|8/1=8
  reg multm_reduce_sa50;  // 9:17|8/1=8
  reg multm_reduce_sa51;  // 9:17|8/1=8
  reg multm_reduce_sa52;  // 9:17|8/1=8
  reg multm_reduce_sa53;  // 9:17|8/1=8
  reg multm_reduce_sa54;  // 9:17|8/1=8
  reg multm_reduce_sa55;  // 9:17|8/1=8
  reg multm_reduce_sa56;  // 9:17|8/1=8
  reg multm_reduce_sa57;  // 9:17|8/1=8
  reg multm_reduce_sa58;  // 9:17|8/1=8
  reg multm_reduce_sa59;  // 9:17|8/1=8
  reg multm_reduce_sa60;  // 9:17|8/1=8
  reg multm_reduce_sa61;  // 9:17|8/1=8
  reg multm_reduce_sa62;  // 9:17|8/1=8
  reg multm_reduce_sa63;  // 9:17|8/1=8
  reg multm_reduce_sa64;  // 9:17|8/1=8
  reg multm_reduce_sa65;  // 9:17|8/1=8
  reg multm_reduce_sa66;  // 9:17|8/1=8
  reg multm_reduce_sa67;  // 9:17|8/1=8
  reg multm_reduce_sa68;  // 9:17|8/1=8
  reg multm_reduce_sa69;  // 9:17|8/1=8
  reg multm_reduce_sa70;  // 9:17|8/1=8
  reg multm_reduce_sa71;  // 9:17|8/1=8
  reg multm_reduce_sa72;  // 9:17|8/1=8
  reg multm_reduce_sa73;  // 9:17|8/1=8
  reg multm_reduce_sa74;  // 9:17|8/1=8
  reg multm_reduce_sa75;  // 9:17|8/1=8
  reg multm_reduce_sa76;  // 9:17|8/1=8
  reg multm_reduce_sa77;  // 9:17|8/1=8
  reg multm_reduce_sa78;  // 9:17|8/1=8
  reg multm_reduce_sa79;  // 9:17|8/1=8
  reg multm_reduce_sa80;  // 9:17|8/1=8
  reg multm_reduce_sa81;  // 9:17|8/1=8
  reg multm_reduce_sa82;  // 9:17|8/1=8
  reg multm_reduce_sa83;  // 9:17|8/1=8
  reg multm_reduce_sa84;  // 9:17|8/1=8
  reg multm_reduce_sa85;  // 9:17|8/1=8
  reg multm_reduce_sa86;  // 9:17|8/1=8
  reg multm_reduce_sa87;  // 9:17|8/1=8
  reg multm_reduce_sa88;  // 9:17|8/1=8
  reg multm_reduce_sa89;  // 9:17|8/1=8
  reg multm_reduce_sa90;  // 9:17|8/1=8
  reg multm_reduce_sa91;  // 9:17|8/1=8
  reg multm_reduce_sa92;  // 9:17|8/1=8
  reg multm_reduce_sa93;  // 9:17|8/1=8
  reg multm_reduce_sa94;  // 9:17|8/1=8
  reg multm_reduce_sa95;  // 9:17|8/1=8
  reg multm_reduce_sa96;  // 9:17|8/1=8
  reg multm_reduce_sa97;  // 9:17|8/1=8
  reg multm_reduce_sa98;  // 9:17|8/1=8
  reg multm_reduce_sa99;  // 9:17|8/1=8
  reg multm_reduce_sa100;  // 9:17|8/1=8
  reg multm_reduce_sa101;  // 9:17|8/1=8
  reg multm_reduce_sa102;  // 9:17|8/1=8
  reg multm_reduce_sa103;  // 9:17|8/1=8
  reg multm_reduce_sa104;  // 9:17|8/1=8
  reg multm_reduce_sa105;  // 9:17|8/1=8
  reg multm_reduce_sa106;  // 9:17|8/1=8
  reg multm_reduce_sa107;  // 9:17|8/1=8
  reg multm_reduce_sa108;  // 9:17|8/1=8
  reg multm_reduce_sa109;  // 9:17|8/1=8
  reg multm_reduce_sa110;  // 9:17|8/1=8
  reg multm_reduce_sa111;  // 9:17|8/1=8
  reg multm_reduce_sa112;  // 9:17|8/1=8
  reg multm_reduce_sa113;  // 9:17|8/1=8
  reg multm_reduce_sa114;  // 9:17|8/1=8
  reg multm_reduce_sa115;  // 9:17|8/1=8
  reg multm_reduce_sa116;  // 9:17|8/1=8
  reg multm_reduce_sa117;  // 9:17|8/1=8
  reg multm_reduce_sa118;  // 9:17|8/1=8
  reg multm_reduce_sa119;  // 9:17|8/1=8
  reg multm_reduce_sa120;  // 9:17|8/1=8
  reg multm_reduce_sa121;  // 9:17|8/1=8
  reg multm_reduce_sa122;  // 9:17|8/1=8
  reg multm_reduce_sa123;  // 9:17|8/1=8
  reg multm_reduce_sa124;  // 9:17|8/1=8
  reg multm_reduce_sa125;  // 9:17|8/1=8
  reg multm_reduce_sa126;  // 9:17|8/1=8
  reg multm_reduce_sa127;  // 9:17|8/1=8
  reg multm_reduce_sa128;  // 9:17|8/1=8
  reg multm_reduce_sa129;  // 9:17|8/1=8
  reg multm_reduce_sa130;  // 9:17|8/1=8
  reg multm_reduce_sa131;  // 9:17|8/1=8
  reg multm_reduce_sa132;  // 9:17|8/1=8
  reg multm_reduce_sa133;  // 9:17|8/1=8
  reg multm_reduce_sa134;  // 9:17|8/1=8
  reg multm_reduce_sa135;  // 9:17|8/1=8
  reg multm_reduce_sa136;  // 9:17|8/1=8
  reg multm_reduce_sa137;  // 9:17|8/1=8
  reg multm_reduce_sa138;  // 9:17|8/1=8
  reg multm_reduce_sa139;  // 9:17|8/1=8
  reg multm_reduce_sa140;  // 9:17|8/1=8
  reg multm_reduce_sa141;  // 9:17|8/1=8
  reg multm_reduce_sa142;  // 9:17|8/1=8
  reg multm_reduce_sa143;  // 9:17|8/1=8
  reg multm_reduce_sa144;  // 9:17|8/1=8
  reg multm_reduce_sa145;  // 9:17|8/1=8
  reg multm_reduce_sa146;  // 9:17|8/1=8
  reg multm_reduce_sa147;  // 9:17|8/1=8
  reg multm_reduce_sa148;  // 9:17|8/1=8
  reg multm_reduce_sa149;  // 9:17|8/1=8
  reg multm_reduce_sa150;  // 9:17|8/1=8
  reg multm_reduce_sa151;  // 9:17|8/1=8
  reg multm_reduce_sa152;  // 9:17|8/1=8
  reg multm_reduce_sa153;  // 9:17|8/1=8
  reg multm_reduce_sa154;  // 9:17|8/1=8
  reg multm_reduce_sa155;  // 9:17|8/1=8
  reg multm_reduce_sa156;  // 9:17|8/1=8
  reg multm_reduce_sa157;  // 9:17|8/1=8
  reg multm_reduce_sa158;  // 9:17|8/1=8
  reg multm_reduce_sa159;  // 9:17|8/1=8
  reg multm_reduce_sa160;  // 9:17|8/1=8
  reg multm_reduce_sa161;  // 9:17|8/1=8
  reg multm_reduce_sa162;  // 9:17|8/1=8
  reg multm_reduce_sa163;  // 9:17|8/1=8
  reg multm_reduce_sa164;  // 9:17|8/1=8
  reg multm_reduce_sa165;  // 9:17|8/1=8
  reg multm_reduce_sa166;  // 9:17|8/1=8
  reg multm_reduce_sa167;  // 9:17|8/1=8
  reg multm_reduce_sa168;  // 9:17|8/1=8
  reg multm_reduce_sa169;  // 9:17|8/1=8
  reg multm_reduce_sa170;  // 9:17|8/1=8
  reg multm_reduce_sa171;  // 9:17|8/1=8
  reg multm_reduce_sa172;  // 9:17|8/1=8
  reg multm_reduce_sa173;  // 9:17|8/1=8
  reg multm_reduce_sa174;  // 9:17|8/1=8
  reg multm_reduce_sa175;  // 9:17|8/1=8
  reg multm_reduce_sa176;  // 9:17|8/1=8
  reg multm_reduce_sa177;  // 9:17|8/1=8
  reg multm_reduce_sa178;  // 9:17|8/1=8
  reg multm_reduce_sa179;  // 9:17|8/1=8
  reg multm_reduce_sa180;  // 9:17|8/1=8
  reg multm_reduce_sa181;  // 9:17|8/1=8
  reg multm_reduce_sa182;  // 9:17|8/1=8
  reg multm_reduce_sa183;  // 9:17|8/1=8
  reg multm_reduce_sa184;  // 9:17|6/1=6
  reg multm_reduce_sa185;  // 9:17|5/1=5
  reg multm_reduce_sb0;  // 8:15|6/1=6
  reg multm_reduce_sb1;  // 9:20|6/1=6
  reg multm_reduce_sb2;  // 9:20|6/1=6
  reg multm_reduce_sb3;  // 9:20|6/1=6
  reg multm_reduce_sb4;  // 9:20|6/1=6
  reg multm_reduce_sb5;  // 9:20|6/1=6
  reg multm_reduce_sb6;  // 9:20|6/1=6
  reg multm_reduce_sb7;  // 9:20|6/1=6
  reg multm_reduce_sb8;  // 9:20|6/1=6
  reg multm_reduce_sb9;  // 9:20|6/1=6
  reg multm_reduce_sb10;  // 9:20|6/1=6
  reg multm_reduce_sb11;  // 9:20|6/1=6
  reg multm_reduce_sb12;  // 9:20|6/1=6
  reg multm_reduce_sb13;  // 9:20|6/1=6
  reg multm_reduce_sb14;  // 9:20|6/1=6
  reg multm_reduce_sb15;  // 9:20|6/1=6
  reg multm_reduce_sb16;  // 9:20|6/1=6
  reg multm_reduce_sb17;  // 9:20|6/1=6
  reg multm_reduce_sb18;  // 9:20|6/1=6
  reg multm_reduce_sb19;  // 9:20|6/1=6
  reg multm_reduce_sb20;  // 9:20|6/1=6
  reg multm_reduce_sb21;  // 9:20|6/1=6
  reg multm_reduce_sb22;  // 9:20|6/1=6
  reg multm_reduce_sb23;  // 9:20|6/1=6
  reg multm_reduce_sb24;  // 9:20|6/1=6
  reg multm_reduce_sb25;  // 9:20|6/1=6
  reg multm_reduce_sb26;  // 9:20|6/1=6
  reg multm_reduce_sb27;  // 9:20|6/1=6
  reg multm_reduce_sb28;  // 9:20|6/1=6
  reg multm_reduce_sb29;  // 9:20|6/1=6
  reg multm_reduce_sb30;  // 9:20|6/1=6
  reg multm_reduce_sb31;  // 9:20|6/1=6
  reg multm_reduce_sb32;  // 9:20|6/1=6
  reg multm_reduce_sb33;  // 9:20|6/1=6
  reg multm_reduce_sb34;  // 9:20|6/1=6
  reg multm_reduce_sb35;  // 9:20|6/1=6
  reg multm_reduce_sb36;  // 9:20|6/1=6
  reg multm_reduce_sb37;  // 9:20|6/1=6
  reg multm_reduce_sb38;  // 9:20|6/1=6
  reg multm_reduce_sb39;  // 9:20|6/1=6
  reg multm_reduce_sb40;  // 9:20|6/1=6
  reg multm_reduce_sb41;  // 9:20|6/1=6
  reg multm_reduce_sb42;  // 9:20|6/1=6
  reg multm_reduce_sb43;  // 9:20|6/1=6
  reg multm_reduce_sb44;  // 9:20|6/1=6
  reg multm_reduce_sb45;  // 9:20|6/1=6
  reg multm_reduce_sb46;  // 9:20|6/1=6
  reg multm_reduce_sb47;  // 9:20|6/1=6
  reg multm_reduce_sb48;  // 9:20|6/1=6
  reg multm_reduce_sb49;  // 9:20|6/1=6
  reg multm_reduce_sb50;  // 9:20|6/1=6
  reg multm_reduce_sb51;  // 9:20|6/1=6
  reg multm_reduce_sb52;  // 9:20|6/1=6
  reg multm_reduce_sb53;  // 9:20|6/1=6
  reg multm_reduce_sb54;  // 9:20|6/1=6
  reg multm_reduce_sb55;  // 9:20|6/1=6
  reg multm_reduce_sb56;  // 9:20|6/1=6
  reg multm_reduce_sb57;  // 9:20|6/1=6
  reg multm_reduce_sb58;  // 9:20|6/1=6
  reg multm_reduce_sb59;  // 9:20|6/1=6
  reg multm_reduce_sb60;  // 9:20|6/1=6
  reg multm_reduce_sb61;  // 9:20|6/1=6
  reg multm_reduce_sb62;  // 9:20|6/1=6
  reg multm_reduce_sb63;  // 9:20|6/1=6
  reg multm_reduce_sb64;  // 9:20|6/1=6
  reg multm_reduce_sb65;  // 9:20|6/1=6
  reg multm_reduce_sb66;  // 9:20|6/1=6
  reg multm_reduce_sb67;  // 9:20|6/1=6
  reg multm_reduce_sb68;  // 9:20|6/1=6
  reg multm_reduce_sb69;  // 9:20|6/1=6
  reg multm_reduce_sb70;  // 9:20|6/1=6
  reg multm_reduce_sb71;  // 9:20|6/1=6
  reg multm_reduce_sb72;  // 9:20|6/1=6
  reg multm_reduce_sb73;  // 9:20|6/1=6
  reg multm_reduce_sb74;  // 9:20|6/1=6
  reg multm_reduce_sb75;  // 9:20|6/1=6
  reg multm_reduce_sb76;  // 9:20|6/1=6
  reg multm_reduce_sb77;  // 9:20|6/1=6
  reg multm_reduce_sb78;  // 9:20|6/1=6
  reg multm_reduce_sb79;  // 9:20|6/1=6
  reg multm_reduce_sb80;  // 9:20|6/1=6
  reg multm_reduce_sb81;  // 9:20|6/1=6
  reg multm_reduce_sb82;  // 9:20|6/1=6
  reg multm_reduce_sb83;  // 9:20|6/1=6
  reg multm_reduce_sb84;  // 9:20|6/1=6
  reg multm_reduce_sb85;  // 9:20|6/1=6
  reg multm_reduce_sb86;  // 9:20|6/1=6
  reg multm_reduce_sb87;  // 9:20|6/1=6
  reg multm_reduce_sb88;  // 9:20|6/1=6
  reg multm_reduce_sb89;  // 9:20|6/1=6
  reg multm_reduce_sb90;  // 9:20|6/1=6
  reg multm_reduce_sb91;  // 9:20|6/1=6
  reg multm_reduce_sb92;  // 9:20|6/1=6
  reg multm_reduce_sb93;  // 9:20|6/1=6
  reg multm_reduce_sb94;  // 9:20|6/1=6
  reg multm_reduce_sb95;  // 9:20|6/1=6
  reg multm_reduce_sb96;  // 9:20|6/1=6
  reg multm_reduce_sb97;  // 9:20|6/1=6
  reg multm_reduce_sb98;  // 9:20|6/1=6
  reg multm_reduce_sb99;  // 9:20|6/1=6
  reg multm_reduce_sb100;  // 9:20|6/1=6
  reg multm_reduce_sb101;  // 9:20|6/1=6
  reg multm_reduce_sb102;  // 9:20|6/1=6
  reg multm_reduce_sb103;  // 9:20|6/1=6
  reg multm_reduce_sb104;  // 9:20|6/1=6
  reg multm_reduce_sb105;  // 9:20|6/1=6
  reg multm_reduce_sb106;  // 9:20|6/1=6
  reg multm_reduce_sb107;  // 9:20|6/1=6
  reg multm_reduce_sb108;  // 9:20|6/1=6
  reg multm_reduce_sb109;  // 9:20|6/1=6
  reg multm_reduce_sb110;  // 9:20|6/1=6
  reg multm_reduce_sb111;  // 9:20|6/1=6
  reg multm_reduce_sb112;  // 9:20|6/1=6
  reg multm_reduce_sb113;  // 9:20|6/1=6
  reg multm_reduce_sb114;  // 9:20|6/1=6
  reg multm_reduce_sb115;  // 9:20|6/1=6
  reg multm_reduce_sb116;  // 9:20|6/1=6
  reg multm_reduce_sb117;  // 9:20|6/1=6
  reg multm_reduce_sb118;  // 9:20|6/1=6
  reg multm_reduce_sb119;  // 9:20|6/1=6
  reg multm_reduce_sb120;  // 9:20|6/1=6
  reg multm_reduce_sb121;  // 9:20|6/1=6
  reg multm_reduce_sb122;  // 9:20|6/1=6
  reg multm_reduce_sb123;  // 9:20|6/1=6
  reg multm_reduce_sb124;  // 9:20|6/1=6
  reg multm_reduce_sb125;  // 9:20|6/1=6
  reg multm_reduce_sb126;  // 9:20|6/1=6
  reg multm_reduce_sb127;  // 9:20|6/1=6
  reg multm_reduce_sb128;  // 9:20|6/1=6
  reg multm_reduce_sb129;  // 9:20|6/1=6
  reg multm_reduce_sb130;  // 9:20|6/1=6
  reg multm_reduce_sb131;  // 9:20|6/1=6
  reg multm_reduce_sb132;  // 9:20|6/1=6
  reg multm_reduce_sb133;  // 9:20|6/1=6
  reg multm_reduce_sb134;  // 9:20|6/1=6
  reg multm_reduce_sb135;  // 9:20|6/1=6
  reg multm_reduce_sb136;  // 9:20|6/1=6
  reg multm_reduce_sb137;  // 9:20|6/1=6
  reg multm_reduce_sb138;  // 9:20|6/1=6
  reg multm_reduce_sb139;  // 9:20|6/1=6
  reg multm_reduce_sb140;  // 9:20|6/1=6
  reg multm_reduce_sb141;  // 9:20|6/1=6
  reg multm_reduce_sb142;  // 9:20|6/1=6
  reg multm_reduce_sb143;  // 9:20|6/1=6
  reg multm_reduce_sb144;  // 9:20|6/1=6
  reg multm_reduce_sb145;  // 9:20|6/1=6
  reg multm_reduce_sb146;  // 9:20|6/1=6
  reg multm_reduce_sb147;  // 9:20|6/1=6
  reg multm_reduce_sb148;  // 9:20|6/1=6
  reg multm_reduce_sb149;  // 9:20|6/1=6
  reg multm_reduce_sb150;  // 9:20|6/1=6
  reg multm_reduce_sb151;  // 9:20|6/1=6
  reg multm_reduce_sb152;  // 9:20|6/1=6
  reg multm_reduce_sb153;  // 9:20|6/1=6
  reg multm_reduce_sb154;  // 9:20|6/1=6
  reg multm_reduce_sb155;  // 9:20|6/1=6
  reg multm_reduce_sb156;  // 9:20|6/1=6
  reg multm_reduce_sb157;  // 9:20|6/1=6
  reg multm_reduce_sb158;  // 9:20|6/1=6
  reg multm_reduce_sb159;  // 9:20|6/1=6
  reg multm_reduce_sb160;  // 9:20|6/1=6
  reg multm_reduce_sb161;  // 9:20|6/1=6
  reg multm_reduce_sb162;  // 9:20|6/1=6
  reg multm_reduce_sb163;  // 9:20|6/1=6
  reg multm_reduce_sb164;  // 9:20|6/1=6
  reg multm_reduce_sb165;  // 9:20|6/1=6
  reg multm_reduce_sb166;  // 9:20|6/1=6
  reg multm_reduce_sb167;  // 9:20|6/1=6
  reg multm_reduce_sb168;  // 9:20|6/1=6
  reg multm_reduce_sb169;  // 9:20|6/1=6
  reg multm_reduce_sb170;  // 9:20|6/1=6
  reg multm_reduce_sb171;  // 9:20|6/1=6
  reg multm_reduce_sb172;  // 9:20|6/1=6
  reg multm_reduce_sb173;  // 9:20|6/1=6
  reg multm_reduce_sb174;  // 9:20|5/1=5
  reg multm_reduce_sc0;  // 5:8|5/1=5
  reg multm_reduce_sc1;  // 6:13|6/1=6
  reg multm_reduce_sc2;  // 6:12|6/1=6
  reg multm_reduce_sc3;  // 5:8|6/1=6
  reg multm_reduce_sc4;  // 6:9|6/1=6
  reg multm_reduce_sc5;  // 6:13|6/1=6
  reg multm_reduce_sc6;  // 6:13|6/1=6
  reg multm_reduce_sc7;  // 6:13|6/1=6
  reg multm_reduce_sc8;  // 6:12|6/1=6
  reg multm_reduce_sc9;  // 5:8|6/1=6
  reg multm_reduce_sc10;  // 6:9|7/1=7
  reg multm_reduce_sc11;  // 6:12|8/1=8
  reg multm_reduce_sc12;  // 6:9|8/1=8
  reg multm_reduce_sc13;  // 6:12|8/1=8
  reg multm_reduce_sc14;  // 5:8|8/1=8
  reg multm_reduce_sc15;  // 5:8|8/1=8
  reg multm_reduce_sc16;  // 5:8|8/1=8
  reg multm_reduce_sc17;  // 5:8|8/1=8
  reg multm_reduce_sc18;  // 6:9|8/1=8
  reg multm_reduce_sc19;  // 6:12|8/1=8
  reg multm_reduce_sc20;  // 6:9|8/1=8
  reg multm_reduce_sc21;  // 6:12|8/1=8
  reg multm_reduce_sc22;  // 6:9|8/1=8
  reg multm_reduce_sc23;  // 6:13|8/1=8
  reg multm_reduce_sc24;  // 6:13|8/1=8
  reg multm_reduce_sc25;  // 6:12|8/1=8
  reg multm_reduce_sc26;  // 5:8|8/1=8
  reg multm_reduce_sc27;  // 5:8|8/1=8
  reg multm_reduce_sc28;  // 6:9|8/1=8
  reg multm_reduce_sc29;  // 6:12|8/1=8
  reg multm_reduce_sc30;  // 6:9|8/1=8
  reg multm_reduce_sc31;  // 6:12|8/1=8
  reg multm_reduce_sc32;  // 6:9|8/1=8
  reg multm_reduce_sc33;  // 6:12|8/1=8
  reg multm_reduce_sc34;  // 6:9|8/1=8
  reg multm_reduce_sc35;  // 6:12|8/1=8
  reg multm_reduce_sc36;  // 5:8|8/1=8
  reg multm_reduce_sc37;  // 6:9|8/1=8
  reg multm_reduce_sc38;  // 6:12|8/1=8
  reg multm_reduce_sc39;  // 5:8|8/1=8
  reg multm_reduce_sc40;  // 6:9|8/1=8
  reg multm_reduce_sc41;  // 6:13|8/1=8
  reg multm_reduce_sc42;  // 6:13|8/1=8
  reg multm_reduce_sc43;  // 6:13|8/1=8
  reg multm_reduce_sc44;  // 6:12|8/1=8
  reg multm_reduce_sc45;  // 5:8|8/1=8
  reg multm_reduce_sc46;  // 5:8|8/1=8
  reg multm_reduce_sc47;  // 6:9|8/1=8
  reg multm_reduce_sc48;  // 6:13|8/1=8
  reg multm_reduce_sc49;  // 6:12|8/1=8
  reg multm_reduce_sc50;  // 5:8|8/1=8
  reg multm_reduce_sc51;  // 6:9|8/1=8
  reg multm_reduce_sc52;  // 6:13|8/1=8
  reg multm_reduce_sc53;  // 6:13|8/1=8
  reg multm_reduce_sc54;  // 6:13|8/1=8
  reg multm_reduce_sc55;  // 6:13|8/1=8
  reg multm_reduce_sc56;  // 6:12|8/1=8
  reg multm_reduce_sc57;  // 6:9|8/1=8
  reg multm_reduce_sc58;  // 6:12|8/1=8
  reg multm_reduce_sc59;  // 5:8|8/1=8
  reg multm_reduce_sc60;  // 5:8|8/1=8
  reg multm_reduce_sc61;  // 5:8|8/1=8
  reg multm_reduce_sc62;  // 6:9|8/1=8
  reg multm_reduce_sc63;  // 6:12|8/1=8
  reg multm_reduce_sc64;  // 5:8|8/1=8
  reg multm_reduce_sc65;  // 5:8|8/1=8
  reg multm_reduce_sc66;  // 6:9|8/1=8
  reg multm_reduce_sc67;  // 6:12|8/1=8
  reg multm_reduce_sc68;  // 6:9|8/1=8
  reg multm_reduce_sc69;  // 6:13|8/1=8
  reg multm_reduce_sc70;  // 6:12|8/1=8
  reg multm_reduce_sc71;  // 6:9|8/1=8
  reg multm_reduce_sc72;  // 6:12|8/1=8
  reg multm_reduce_sc73;  // 6:9|8/1=8
  reg multm_reduce_sc74;  // 6:13|8/1=8
  reg multm_reduce_sc75;  // 6:12|8/1=8
  reg multm_reduce_sc76;  // 5:8|8/1=8
  reg multm_reduce_sc77;  // 5:8|8/1=8
  reg multm_reduce_sc78;  // 5:8|8/1=8
  reg multm_reduce_sc79;  // 6:9|8/1=8
  reg multm_reduce_sc80;  // 6:13|8/1=8
  reg multm_reduce_sc81;  // 6:12|8/1=8
  reg multm_reduce_sc82;  // 6:9|8/1=8
  reg multm_reduce_sc83;  // 6:12|8/1=8
  reg multm_reduce_sc84;  // 5:8|8/1=8
  reg multm_reduce_sc85;  // 5:8|8/1=8
  reg multm_reduce_sc86;  // 6:9|8/1=8
  reg multm_reduce_sc87;  // 6:12|8/1=8
  reg multm_reduce_sc88;  // 6:9|8/1=8
  reg multm_reduce_sc89;  // 6:12|8/1=8
  reg multm_reduce_sc90;  // 6:9|8/1=8
  reg multm_reduce_sc91;  // 6:13|8/1=8
  reg multm_reduce_sc92;  // 6:12|8/1=8
  reg multm_reduce_sc93;  // 5:8|8/1=8
  reg multm_reduce_sc94;  // 5:8|8/1=8
  reg multm_reduce_sc95;  // 5:8|8/1=8
  reg multm_reduce_sc96;  // 6:9|8/1=8
  reg multm_reduce_sc97;  // 6:12|8/1=8
  reg multm_reduce_sc98;  // 5:8|8/1=8
  reg multm_reduce_sc99;  // 6:9|8/1=8
  reg multm_reduce_sc100;  // 6:13|8/1=8
  reg multm_reduce_sc101;  // 6:13|8/1=8
  reg multm_reduce_sc102;  // 6:13|8/1=8
  reg multm_reduce_sc103;  // 6:12|8/1=8
  reg multm_reduce_sc104;  // 6:9|8/1=8
  reg multm_reduce_sc105;  // 6:13|8/1=8
  reg multm_reduce_sc106;  // 6:12|8/1=8
  reg multm_reduce_sc107;  // 6:9|8/1=8
  reg multm_reduce_sc108;  // 6:13|8/1=8
  reg multm_reduce_sc109;  // 6:13|8/1=8
  reg multm_reduce_sc110;  // 6:13|8/1=8
  reg multm_reduce_sc111;  // 6:12|8/1=8
  reg multm_reduce_sc112;  // 6:9|8/1=8
  reg multm_reduce_sc113;  // 6:12|8/1=8
  reg multm_reduce_sc114;  // 6:9|8/1=8
  reg multm_reduce_sc115;  // 6:12|8/1=8
  reg multm_reduce_sc116;  // 5:8|8/1=8
  reg multm_reduce_sc117;  // 6:9|8/1=8
  reg multm_reduce_sc118;  // 6:13|8/1=8
  reg multm_reduce_sc119;  // 6:13|8/1=8
  reg multm_reduce_sc120;  // 6:13|8/1=8
  reg multm_reduce_sc121;  // 6:13|8/1=8
  reg multm_reduce_sc122;  // 6:13|8/1=8
  reg multm_reduce_sc123;  // 6:13|8/1=8
  reg multm_reduce_sc124;  // 6:12|8/1=8
  reg multm_reduce_sc125;  // 5:8|8/1=8
  reg multm_reduce_sc126;  // 5:8|8/1=8
  reg multm_reduce_sc127;  // 5:8|8/1=8
  reg multm_reduce_sc128;  // 6:9|8/1=8
  reg multm_reduce_sc129;  // 6:12|8/1=8
  reg multm_reduce_sc130;  // 6:9|8/1=8
  reg multm_reduce_sc131;  // 6:12|8/1=8
  reg multm_reduce_sc132;  // 6:9|8/1=8
  reg multm_reduce_sc133;  // 6:12|8/1=8
  reg multm_reduce_sc134;  // 5:8|8/1=8
  reg multm_reduce_sc135;  // 6:9|8/1=8
  reg multm_reduce_sc136;  // 6:13|8/1=8
  reg multm_reduce_sc137;  // 6:12|8/1=8
  reg multm_reduce_sc138;  // 5:8|8/1=8
  reg multm_reduce_sc139;  // 5:8|8/1=8
  reg multm_reduce_sc140;  // 6:9|8/1=8
  reg multm_reduce_sc141;  // 6:13|8/1=8
  reg multm_reduce_sc142;  // 6:13|8/1=8
  reg multm_reduce_sc143;  // 6:13|8/1=8
  reg multm_reduce_sc144;  // 6:13|8/1=8
  reg multm_reduce_sc145;  // 6:12|8/1=8
  reg multm_reduce_sc146;  // 5:8|8/1=8
  reg multm_reduce_sc147;  // 6:9|8/1=8
  reg multm_reduce_sc148;  // 6:12|8/1=8
  reg multm_reduce_sc149;  // 5:8|8/1=8
  reg multm_reduce_sc150;  // 6:9|8/1=8
  reg multm_reduce_sc151;  // 6:13|8/1=8
  reg multm_reduce_sc152;  // 6:13|8/1=8
  reg multm_reduce_sc153;  // 6:13|8/1=8
  reg multm_reduce_sc154;  // 6:12|8/1=8
  reg multm_reduce_sc155;  // 6:9|8/1=8
  reg multm_reduce_sc156;  // 6:13|8/1=8
  reg multm_reduce_sc157;  // 6:13|8/1=8
  reg multm_reduce_sc158;  // 6:13|8/1=8
  reg multm_reduce_sc159;  // 6:13|8/1=8
  reg multm_reduce_sc160;  // 6:13|8/1=8
  reg multm_reduce_sc161;  // 6:12|8/1=8
  reg multm_reduce_sc162;  // 6:9|8/1=8
  reg multm_reduce_sc163;  // 6:12|8/1=8
  reg multm_reduce_sc164;  // 5:8|8/1=8
  reg multm_reduce_sc165;  // 5:8|8/1=8
  reg multm_reduce_sc166;  // 6:9|8/1=8
  reg multm_reduce_sc167;  // 6:12|8/1=8
  reg multm_reduce_sc168;  // 5:8|8/1=8
  reg multm_reduce_sc169;  // 5:8|8/1=8
  reg multm_reduce_sc170;  // 5:8|8/1=8
  reg multm_reduce_sc171;  // 6:9|8/1=8
  reg multm_reduce_sc172;  // 6:13|8/1=8
  reg multm_reduce_sc173;  // 6:13|8/1=8
  reg multm_reduce_sc174;  // 6:13|8/1=8
  reg multm_reduce_sc175;  // 6:13|8/1=8
  reg multm_reduce_sc176;  // 6:12|8/1=8
  reg multm_reduce_sc177;  // 5:8|8/1=8
  reg multm_reduce_sc178;  // 5:8|8/1=8
  reg multm_reduce_sc179;  // 6:9|8/1=8
  reg multm_reduce_sc180;  // 6:12|8/1=8
  reg multm_reduce_sc181;  // 6:9|8/1=8
  reg multm_reduce_sc182;  // 5:11|8/1=8
  reg multm_reduce_sd0;  // 4:5|3/1=3
  reg multm_reduce_sd1;  // 5:8|6/1=6
  reg multm_reduce_sd2;  // 6:13|6/1=6
  reg multm_reduce_sd3;  // 6:12|6/1=6
  reg multm_reduce_sd4;  // 5:8|6/1=6
  reg multm_reduce_sd5;  // 6:9|6/1=6
  reg multm_reduce_sd6;  // 6:13|6/1=6
  reg multm_reduce_sd7;  // 6:13|6/1=6
  reg multm_reduce_sd8;  // 6:13|6/1=6
  reg multm_reduce_sd9;  // 6:12|6/1=6
  reg multm_reduce_sd10;  // 5:8|7/1=7
  reg multm_reduce_sd11;  // 6:9|8/1=8
  reg multm_reduce_sd12;  // 6:12|8/1=8
  reg multm_reduce_sd13;  // 6:9|8/1=8
  reg multm_reduce_sd14;  // 6:12|8/1=8
  reg multm_reduce_sd15;  // 5:8|8/1=8
  reg multm_reduce_sd16;  // 5:8|8/1=8
  reg multm_reduce_sd17;  // 5:8|8/1=8
  reg multm_reduce_sd18;  // 5:8|8/1=8
  reg multm_reduce_sd19;  // 6:9|8/1=8
  reg multm_reduce_sd20;  // 6:12|8/1=8
  reg multm_reduce_sd21;  // 6:9|8/1=8
  reg multm_reduce_sd22;  // 6:12|8/1=8
  reg multm_reduce_sd23;  // 6:9|8/1=8
  reg multm_reduce_sd24;  // 6:13|8/1=8
  reg multm_reduce_sd25;  // 6:13|8/1=8
  reg multm_reduce_sd26;  // 6:12|8/1=8
  reg multm_reduce_sd27;  // 5:8|8/1=8
  reg multm_reduce_sd28;  // 5:8|8/1=8
  reg multm_reduce_sd29;  // 6:9|8/1=8
  reg multm_reduce_sd30;  // 6:12|8/1=8
  reg multm_reduce_sd31;  // 6:9|8/1=8
  reg multm_reduce_sd32;  // 6:12|8/1=8
  reg multm_reduce_sd33;  // 6:9|8/1=8
  reg multm_reduce_sd34;  // 6:12|8/1=8
  reg multm_reduce_sd35;  // 6:9|8/1=8
  reg multm_reduce_sd36;  // 6:12|8/1=8
  reg multm_reduce_sd37;  // 5:8|8/1=8
  reg multm_reduce_sd38;  // 6:9|8/1=8
  reg multm_reduce_sd39;  // 6:12|8/1=8
  reg multm_reduce_sd40;  // 5:8|8/1=8
  reg multm_reduce_sd41;  // 6:9|8/1=8
  reg multm_reduce_sd42;  // 6:13|8/1=8
  reg multm_reduce_sd43;  // 6:13|8/1=8
  reg multm_reduce_sd44;  // 6:13|8/1=8
  reg multm_reduce_sd45;  // 6:12|8/1=8
  reg multm_reduce_sd46;  // 5:8|8/1=8
  reg multm_reduce_sd47;  // 5:8|8/1=8
  reg multm_reduce_sd48;  // 6:9|8/1=8
  reg multm_reduce_sd49;  // 6:13|8/1=8
  reg multm_reduce_sd50;  // 6:12|8/1=8
  reg multm_reduce_sd51;  // 5:8|8/1=8
  reg multm_reduce_sd52;  // 6:9|8/1=8
  reg multm_reduce_sd53;  // 6:13|8/1=8
  reg multm_reduce_sd54;  // 6:13|8/1=8
  reg multm_reduce_sd55;  // 6:13|8/1=8
  reg multm_reduce_sd56;  // 6:13|8/1=8
  reg multm_reduce_sd57;  // 6:12|8/1=8
  reg multm_reduce_sd58;  // 6:9|8/1=8
  reg multm_reduce_sd59;  // 6:12|8/1=8
  reg multm_reduce_sd60;  // 5:8|8/1=8
  reg multm_reduce_sd61;  // 5:8|8/1=8
  reg multm_reduce_sd62;  // 5:8|8/1=8
  reg multm_reduce_sd63;  // 6:9|8/1=8
  reg multm_reduce_sd64;  // 6:12|8/1=8
  reg multm_reduce_sd65;  // 5:8|8/1=8
  reg multm_reduce_sd66;  // 5:8|8/1=8
  reg multm_reduce_sd67;  // 6:9|8/1=8
  reg multm_reduce_sd68;  // 6:12|8/1=8
  reg multm_reduce_sd69;  // 6:9|8/1=8
  reg multm_reduce_sd70;  // 6:13|8/1=8
  reg multm_reduce_sd71;  // 6:12|8/1=8
  reg multm_reduce_sd72;  // 6:9|8/1=8
  reg multm_reduce_sd73;  // 6:12|8/1=8
  reg multm_reduce_sd74;  // 6:9|8/1=8
  reg multm_reduce_sd75;  // 6:13|8/1=8
  reg multm_reduce_sd76;  // 6:12|8/1=8
  reg multm_reduce_sd77;  // 5:8|8/1=8
  reg multm_reduce_sd78;  // 5:8|8/1=8
  reg multm_reduce_sd79;  // 5:8|8/1=8
  reg multm_reduce_sd80;  // 6:9|8/1=8
  reg multm_reduce_sd81;  // 6:13|8/1=8
  reg multm_reduce_sd82;  // 6:12|8/1=8
  reg multm_reduce_sd83;  // 6:9|8/1=8
  reg multm_reduce_sd84;  // 6:12|8/1=8
  reg multm_reduce_sd85;  // 5:8|8/1=8
  reg multm_reduce_sd86;  // 5:8|8/1=8
  reg multm_reduce_sd87;  // 6:9|8/1=8
  reg multm_reduce_sd88;  // 6:12|8/1=8
  reg multm_reduce_sd89;  // 6:9|8/1=8
  reg multm_reduce_sd90;  // 6:12|8/1=8
  reg multm_reduce_sd91;  // 6:9|8/1=8
  reg multm_reduce_sd92;  // 6:13|8/1=8
  reg multm_reduce_sd93;  // 6:12|8/1=8
  reg multm_reduce_sd94;  // 5:8|8/1=8
  reg multm_reduce_sd95;  // 5:8|8/1=8
  reg multm_reduce_sd96;  // 5:8|8/1=8
  reg multm_reduce_sd97;  // 6:9|8/1=8
  reg multm_reduce_sd98;  // 6:12|8/1=8
  reg multm_reduce_sd99;  // 5:8|8/1=8
  reg multm_reduce_sd100;  // 6:9|8/1=8
  reg multm_reduce_sd101;  // 6:13|8/1=8
  reg multm_reduce_sd102;  // 6:13|8/1=8
  reg multm_reduce_sd103;  // 6:13|8/1=8
  reg multm_reduce_sd104;  // 6:12|8/1=8
  reg multm_reduce_sd105;  // 6:9|8/1=8
  reg multm_reduce_sd106;  // 6:13|8/1=8
  reg multm_reduce_sd107;  // 6:12|8/1=8
  reg multm_reduce_sd108;  // 6:9|8/1=8
  reg multm_reduce_sd109;  // 6:13|8/1=8
  reg multm_reduce_sd110;  // 6:13|8/1=8
  reg multm_reduce_sd111;  // 6:13|8/1=8
  reg multm_reduce_sd112;  // 6:12|8/1=8
  reg multm_reduce_sd113;  // 6:9|8/1=8
  reg multm_reduce_sd114;  // 6:12|8/1=8
  reg multm_reduce_sd115;  // 6:9|8/1=8
  reg multm_reduce_sd116;  // 6:12|8/1=8
  reg multm_reduce_sd117;  // 5:8|8/1=8
  reg multm_reduce_sd118;  // 6:9|8/1=8
  reg multm_reduce_sd119;  // 6:13|8/1=8
  reg multm_reduce_sd120;  // 6:13|8/1=8
  reg multm_reduce_sd121;  // 6:13|8/1=8
  reg multm_reduce_sd122;  // 6:13|8/1=8
  reg multm_reduce_sd123;  // 6:13|8/1=8
  reg multm_reduce_sd124;  // 6:13|8/1=8
  reg multm_reduce_sd125;  // 6:12|8/1=8
  reg multm_reduce_sd126;  // 5:8|8/1=8
  reg multm_reduce_sd127;  // 5:8|8/1=8
  reg multm_reduce_sd128;  // 5:8|8/1=8
  reg multm_reduce_sd129;  // 6:9|8/1=8
  reg multm_reduce_sd130;  // 6:12|8/1=8
  reg multm_reduce_sd131;  // 6:9|8/1=8
  reg multm_reduce_sd132;  // 6:12|8/1=8
  reg multm_reduce_sd133;  // 6:9|8/1=8
  reg multm_reduce_sd134;  // 6:12|8/1=8
  reg multm_reduce_sd135;  // 5:8|8/1=8
  reg multm_reduce_sd136;  // 6:9|8/1=8
  reg multm_reduce_sd137;  // 6:13|8/1=8
  reg multm_reduce_sd138;  // 6:12|8/1=8
  reg multm_reduce_sd139;  // 5:8|8/1=8
  reg multm_reduce_sd140;  // 5:8|8/1=8
  reg multm_reduce_sd141;  // 6:9|8/1=8
  reg multm_reduce_sd142;  // 6:13|8/1=8
  reg multm_reduce_sd143;  // 6:13|8/1=8
  reg multm_reduce_sd144;  // 6:13|8/1=8
  reg multm_reduce_sd145;  // 6:13|8/1=8
  reg multm_reduce_sd146;  // 6:12|8/1=8
  reg multm_reduce_sd147;  // 5:8|8/1=8
  reg multm_reduce_sd148;  // 6:9|8/1=8
  reg multm_reduce_sd149;  // 6:12|8/1=8
  reg multm_reduce_sd150;  // 5:8|8/1=8
  reg multm_reduce_sd151;  // 6:9|8/1=8
  reg multm_reduce_sd152;  // 6:13|8/1=8
  reg multm_reduce_sd153;  // 6:13|8/1=8
  reg multm_reduce_sd154;  // 6:13|8/1=8
  reg multm_reduce_sd155;  // 6:12|8/1=8
  reg multm_reduce_sd156;  // 6:9|8/1=8
  reg multm_reduce_sd157;  // 6:13|8/1=8
  reg multm_reduce_sd158;  // 6:13|8/1=8
  reg multm_reduce_sd159;  // 6:13|8/1=8
  reg multm_reduce_sd160;  // 6:13|8/1=8
  reg multm_reduce_sd161;  // 6:13|8/1=8
  reg multm_reduce_sd162;  // 6:12|8/1=8
  reg multm_reduce_sd163;  // 6:9|8/1=8
  reg multm_reduce_sd164;  // 6:12|8/1=8
  reg multm_reduce_sd165;  // 5:8|8/1=8
  reg multm_reduce_sd166;  // 5:8|8/1=8
  reg multm_reduce_sd167;  // 6:9|8/1=8
  reg multm_reduce_sd168;  // 6:12|8/1=8
  reg multm_reduce_sd169;  // 5:8|8/1=8
  reg multm_reduce_sd170;  // 5:8|8/1=8
  reg multm_reduce_sd171;  // 5:8|8/1=8
  reg multm_reduce_sd172;  // 6:9|8/1=8
  reg multm_reduce_sd173;  // 6:13|8/1=8
  reg multm_reduce_sd174;  // 6:13|8/1=8
  reg multm_reduce_sd175;  // 6:13|8/1=8
  reg multm_reduce_sd176;  // 6:13|8/1=8
  reg multm_reduce_sd177;  // 6:12|8/1=8
  reg multm_reduce_sd178;  // 5:8|8/1=8
  reg multm_reduce_sd179;  // 5:8|8/1=8
  reg multm_reduce_sd180;  // 6:9|8/1=8
  reg multm_reduce_sd181;  // 6:12|8/1=8
  reg multm_reduce_sd182;  // 6:9|8/1=8
  reg multm_reduce_sd183;  // 5:14|6/1=6
  reg pipe0_x1;  // 1:0|1/1=1
  reg pipe0_x2;  // 1:0|1/1=1
  reg pipe0_x3;  // 1:0|1/1=1
  reg pipe0_x4;  // 1:0|1/1=1
  reg pipe0_x5;  // 1:0|1/1=1
  reg pipe0_x6;  // 1:0|1/1=1
  reg pipe0_x7;  // 1:0|1/1=3
  reg pipe0_x8;  // 1:0|1/3=5
  reg pipe0_x9;  // 1:0|1/15=5
  reg pipe1_x1;  // 1:0|1/1=1
  reg pipe1_x2;  // 1:0|1/1=1
  reg pipe1_x3;  // 1:0|1/1=1
  reg pipe1_x4;  // 1:0|1/1=1
  reg pipe1_x5;  // 1:0|1/1=1
  reg pipe1_x6;  // 1:0|1/1=1
  reg pipe1_x7;  // 1:0|1/1=3
  reg pipe1_x8;  // 1:0|1/3=4
  reg pipe1_x9;  // 1:0|1/14=5
  reg sa;  // 6:9|3/1=3
  reg sad;  // 1:0|370/81=5
  reg sadd;  // 1:0|409/74=5
  reg sb;  // 9:14|3/1=3
  reg sbd;  // 1:0|370/72=5
  reg sbdd;  // 1:0|22/4=5
  reg yc0_o;  // 6:3|5/1=5
  reg yc1_o;  // 7:7|5/1=5
  reg yc2_o;  // 6:3|5/1=5
  reg yc3_o;  // 7:7|5/1=5
  reg yc4_o;  // 8:9|5/1=5
  reg yc5_o;  // 8:9|5/1=5
  reg yc6_o;  // 8:8|5/1=5
  reg yc7_o;  // 6:3|5/1=5
  reg yc8_o;  // 6:3|5/1=5
  reg yc9_o;  // 7:7|5/1=5
  reg yc10_o;  // 8:9|5/1=5
  reg yc11_o;  // 8:9|5/1=5
  reg yc12_o;  // 8:9|5/1=5
  reg yc13_o;  // 8:9|5/1=5
  reg yc14_o;  // 8:9|5/1=5
  reg yc15_o;  // 8:8|5/1=5
  reg yc16_o;  // 8:8|5/1=5
  reg yc17_o;  // 8:8|5/1=5
  reg yc18_o;  // 8:8|5/1=5
  reg yc19_o;  // 8:9|5/1=5
  reg yc20_o;  // 8:9|5/1=5
  reg yc21_o;  // 8:9|5/1=5
  reg yc22_o;  // 8:9|5/1=5
  reg yc23_o;  // 8:9|5/1=5
  reg yc24_o;  // 8:8|5/1=5
  reg yc25_o;  // 6:3|5/1=5
  reg yc26_o;  // 7:7|5/1=5
  reg yc27_o;  // 8:9|5/1=5
  reg yc28_o;  // 8:8|5/1=5
  reg yc29_o;  // 8:9|5/1=5
  reg yc30_o;  // 8:9|5/1=5
  reg yc31_o;  // 8:9|5/1=5
  reg yc32_o;  // 8:9|5/1=5
  reg yc33_o;  // 8:9|5/1=5
  reg yc34_o;  // 8:9|5/1=5
  reg yc35_o;  // 8:9|5/1=5
  reg yc36_o;  // 8:9|5/1=5
  reg yc37_o;  // 8:8|5/1=5
  reg yc38_o;  // 8:9|5/1=5
  reg yc39_o;  // 8:9|5/1=5
  reg yc40_o;  // 8:8|5/1=5
  reg yc41_o;  // 8:9|5/1=5
  reg yc42_o;  // 8:8|5/1=5
  reg yc43_o;  // 6:3|5/1=5
  reg yc44_o;  // 6:3|5/1=5
  reg yc45_o;  // 7:7|5/1=5
  reg yc46_o;  // 8:9|5/1=5
  reg yc47_o;  // 8:8|5/1=5
  reg yc48_o;  // 8:9|5/1=5
  reg yc49_o;  // 8:8|5/1=5
  reg yc50_o;  // 7:7|5/1=5
  reg yc51_o;  // 8:9|5/1=5
  reg yc52_o;  // 8:9|5/1=5
  reg yc53_o;  // 8:8|5/1=5
  reg yc54_o;  // 6:3|5/1=5
  reg yc55_o;  // 6:3|5/1=5
  reg yc56_o;  // 6:3|5/1=5
  reg yc57_o;  // 7:7|5/1=5
  reg yc58_o;  // 7:7|5/1=5
  reg yc59_o;  // 7:7|5/1=5
  reg yc60_o;  // 8:9|5/1=5
  reg yc61_o;  // 8:8|5/1=5
  reg yc62_o;  // 8:8|5/1=5
  reg yc63_o;  // 8:9|5/1=5
  reg yc64_o;  // 8:9|5/1=5
  reg yc65_o;  // 8:8|5/1=5
  reg yc66_o;  // 8:8|5/1=5
  reg yc67_o;  // 8:9|5/1=5
  reg yc68_o;  // 8:9|5/1=5
  reg yc69_o;  // 8:9|5/1=5
  reg yc70_o;  // 8:8|5/1=5
  reg yc71_o;  // 7:7|5/1=5
  reg yc72_o;  // 7:7|5/1=5
  reg yc73_o;  // 7:7|5/1=5
  reg yc74_o;  // 7:7|5/1=5
  reg yc75_o;  // 6:3|5/1=5
  reg yc76_o;  // 7:7|5/1=5
  reg yc77_o;  // 8:9|5/1=5
  reg yc78_o;  // 8:8|5/1=5
  reg yc79_o;  // 8:8|5/1=5
  reg yc80_o;  // 8:9|5/1=5
  reg yc81_o;  // 8:8|5/1=5
  reg yc82_o;  // 7:7|5/1=5
  reg yc83_o;  // 7:7|5/1=5
  reg yc84_o;  // 7:7|5/1=5
  reg yc85_o;  // 8:9|5/1=5
  reg yc86_o;  // 8:8|5/1=5
  reg yc87_o;  // 8:9|5/1=5
  reg yc88_o;  // 8:9|5/1=5
  reg yc89_o;  // 8:9|5/1=5
  reg yc90_o;  // 8:9|5/1=5
  reg yc91_o;  // 8:9|5/1=5
  reg yc92_o;  // 8:8|5/1=5
  reg yc93_o;  // 7:7|5/1=5
  reg yc94_o;  // 8:9|5/1=5
  reg yc95_o;  // 8:8|5/1=5
  reg yc96_o;  // 8:8|5/1=5
  reg yc97_o;  // 8:9|5/1=5
  reg yc98_o;  // 8:9|5/1=5
  reg yc99_o;  // 8:8|5/1=5
  reg yc100_o;  // 8:9|5/1=5
  reg yc101_o;  // 8:8|5/1=5
  reg yc102_o;  // 6:3|5/1=5
  reg yc103_o;  // 6:3|5/1=5
  reg yc104_o;  // 7:7|5/1=5
  reg yc105_o;  // 7:7|5/1=5
  reg yc106_o;  // 6:3|5/1=5
  reg yc107_o;  // 7:7|5/1=5
  reg yc108_o;  // 7:7|5/1=5
  reg yc109_o;  // 6:3|5/1=5
  reg yc110_o;  // 6:3|5/1=5
  reg yc111_o;  // 6:3|5/1=5
  reg yc112_o;  // 7:7|5/1=5
  reg yc113_o;  // 7:7|5/1=5
  reg yc114_o;  // 7:7|5/1=5
  reg yc115_o;  // 7:7|5/1=5
  reg yc116_o;  // 7:7|5/1=5
  reg yc117_o;  // 8:9|5/1=5
  reg yc118_o;  // 8:9|5/1=5
  reg yc119_o;  // 8:8|5/1=5
  reg yc120_o;  // 6:3|5/1=5
  reg yc121_o;  // 6:3|5/1=5
  reg yc122_o;  // 6:3|5/1=5
  reg yc123_o;  // 6:3|5/1=5
  reg yc124_o;  // 6:3|5/1=5
  reg yc125_o;  // 7:7|5/1=5
  reg yc126_o;  // 8:9|5/1=5
  reg yc127_o;  // 8:8|5/1=5
  reg yc128_o;  // 8:8|5/1=5
  reg yc129_o;  // 8:9|5/1=5
  reg yc130_o;  // 8:9|5/1=5
  reg yc131_o;  // 8:9|5/1=5
  reg yc132_o;  // 8:9|5/1=5
  reg yc133_o;  // 8:9|5/1=5
  reg yc134_o;  // 8:9|5/1=5
  reg yc135_o;  // 8:8|5/1=5
  reg yc136_o;  // 8:9|5/1=5
  reg yc137_o;  // 8:8|5/1=5
  reg yc138_o;  // 7:7|5/1=5
  reg yc139_o;  // 8:9|5/1=5
  reg yc140_o;  // 8:8|5/1=5
  reg yc141_o;  // 8:9|5/1=5
  reg yc142_o;  // 8:8|5/1=5
  reg yc143_o;  // 6:3|5/1=5
  reg yc144_o;  // 6:3|5/1=5
  reg yc145_o;  // 6:3|5/1=5
  reg yc146_o;  // 7:7|5/1=5
  reg yc147_o;  // 8:9|5/1=5
  reg yc148_o;  // 8:9|5/1=5
  reg yc149_o;  // 8:9|5/1=5
  reg yc150_o;  // 8:8|5/1=5
  reg yc151_o;  // 8:9|5/1=5
  reg yc152_o;  // 8:8|5/1=5
  reg yc153_o;  // 6:3|5/1=5
  reg yc154_o;  // 6:3|5/1=5
  reg yc155_o;  // 7:7|5/1=5
  reg yc156_o;  // 7:7|5/1=5
  reg yc157_o;  // 6:3|5/1=5
  reg yc158_o;  // 6:3|5/1=5
  reg yc159_o;  // 6:3|5/1=5
  reg yc160_o;  // 6:3|5/1=5
  reg yc161_o;  // 6:3|5/1=5
  reg yc162_o;  // 7:7|5/1=5
  reg yc163_o;  // 7:7|5/1=5
  reg yc164_o;  // 7:7|5/1=5
  reg yc165_o;  // 8:9|5/1=5
  reg yc166_o;  // 8:8|5/1=5
  reg yc167_o;  // 8:9|5/1=5
  reg yc168_o;  // 8:9|5/1=5
  reg yc169_o;  // 8:8|5/1=5
  reg yc170_o;  // 8:8|5/1=5
  reg yc171_o;  // 8:8|5/1=5
  reg yc172_o;  // 8:9|5/1=5
  reg yc173_o;  // 8:8|5/1=5
  reg yc174_o;  // 6:3|5/1=5
  reg yc175_o;  // 6:3|5/1=5
  reg yc176_o;  // 6:3|5/1=5
  reg yc177_o;  // 7:7|5/1=5
  reg yc178_o;  // 8:9|5/1=5
  reg yc179_o;  // 8:8|5/1=5
  reg yc180_o;  // 8:9|5/1=5
  reg yc181_o;  // 8:9|5/1=5
  reg yc182_o;  // 8:9|5/1=5
  reg yc183_o;  // 8:8|5/1=5
  reg ys0_o;  // 6:3|6/1=6
  reg ys1_o;  // 7:4|7/1=7
  reg ys2_o;  // 6:3|7/1=7
  reg ys3_o;  // 7:4|7/1=7
  reg ys4_o;  // 8:6|7/1=7
  reg ys5_o;  // 8:6|7/1=7
  reg ys6_o;  // 8:5|7/1=7
  reg ys7_o;  // 6:3|7/1=7
  reg ys8_o;  // 6:3|7/1=7
  reg ys9_o;  // 7:4|7/1=7
  reg ys10_o;  // 8:6|7/1=7
  reg ys11_o;  // 8:6|7/1=7
  reg ys12_o;  // 8:6|7/1=7
  reg ys13_o;  // 8:6|7/1=7
  reg ys14_o;  // 8:6|7/1=7
  reg ys15_o;  // 8:5|7/1=7
  reg ys16_o;  // 8:5|7/1=7
  reg ys17_o;  // 8:5|7/1=7
  reg ys18_o;  // 8:5|7/1=7
  reg ys19_o;  // 8:6|7/1=7
  reg ys20_o;  // 8:6|7/1=7
  reg ys21_o;  // 8:6|7/1=7
  reg ys22_o;  // 8:6|7/1=7
  reg ys23_o;  // 8:6|7/1=7
  reg ys24_o;  // 8:5|7/1=7
  reg ys25_o;  // 6:3|7/1=7
  reg ys26_o;  // 7:4|7/1=7
  reg ys27_o;  // 8:6|7/1=7
  reg ys28_o;  // 8:5|7/1=7
  reg ys29_o;  // 8:6|7/1=7
  reg ys30_o;  // 8:6|7/1=7
  reg ys31_o;  // 8:6|7/1=7
  reg ys32_o;  // 8:6|7/1=7
  reg ys33_o;  // 8:6|7/1=7
  reg ys34_o;  // 8:6|7/1=7
  reg ys35_o;  // 8:6|7/1=7
  reg ys36_o;  // 8:6|7/1=7
  reg ys37_o;  // 8:5|7/1=7
  reg ys38_o;  // 8:6|7/1=7
  reg ys39_o;  // 8:6|7/1=7
  reg ys40_o;  // 8:5|7/1=7
  reg ys41_o;  // 8:6|7/1=7
  reg ys42_o;  // 8:5|7/1=7
  reg ys43_o;  // 6:3|7/1=7
  reg ys44_o;  // 6:3|7/1=7
  reg ys45_o;  // 7:4|7/1=7
  reg ys46_o;  // 8:6|7/1=7
  reg ys47_o;  // 8:5|7/1=7
  reg ys48_o;  // 8:6|7/1=7
  reg ys49_o;  // 8:5|7/1=7
  reg ys50_o;  // 7:4|7/1=7
  reg ys51_o;  // 8:6|7/1=7
  reg ys52_o;  // 8:6|7/1=7
  reg ys53_o;  // 8:5|7/1=7
  reg ys54_o;  // 6:3|7/1=7
  reg ys55_o;  // 6:3|7/1=7
  reg ys56_o;  // 6:3|7/1=7
  reg ys57_o;  // 7:4|7/1=7
  reg ys58_o;  // 7:4|7/1=7
  reg ys59_o;  // 7:4|7/1=7
  reg ys60_o;  // 8:6|7/1=7
  reg ys61_o;  // 8:5|7/1=7
  reg ys62_o;  // 8:5|7/1=7
  reg ys63_o;  // 8:6|7/1=7
  reg ys64_o;  // 8:6|7/1=7
  reg ys65_o;  // 8:5|7/1=7
  reg ys66_o;  // 8:5|7/1=7
  reg ys67_o;  // 8:6|7/1=7
  reg ys68_o;  // 8:6|7/1=7
  reg ys69_o;  // 8:6|7/1=7
  reg ys70_o;  // 8:5|7/1=7
  reg ys71_o;  // 7:4|7/1=7
  reg ys72_o;  // 7:4|7/1=7
  reg ys73_o;  // 7:4|7/1=7
  reg ys74_o;  // 7:4|7/1=7
  reg ys75_o;  // 6:3|7/1=7
  reg ys76_o;  // 7:4|7/1=7
  reg ys77_o;  // 8:6|7/1=7
  reg ys78_o;  // 8:5|7/1=7
  reg ys79_o;  // 8:5|7/1=7
  reg ys80_o;  // 8:6|7/1=7
  reg ys81_o;  // 8:5|7/1=7
  reg ys82_o;  // 7:4|7/1=7
  reg ys83_o;  // 7:4|7/1=7
  reg ys84_o;  // 7:4|7/1=7
  reg ys85_o;  // 8:6|7/1=7
  reg ys86_o;  // 8:5|7/1=7
  reg ys87_o;  // 8:6|7/1=7
  reg ys88_o;  // 8:6|7/1=7
  reg ys89_o;  // 8:6|7/1=7
  reg ys90_o;  // 8:6|7/1=7
  reg ys91_o;  // 8:6|7/1=7
  reg ys92_o;  // 8:5|7/1=7
  reg ys93_o;  // 7:4|7/1=7
  reg ys94_o;  // 8:6|7/1=7
  reg ys95_o;  // 8:5|7/1=7
  reg ys96_o;  // 8:5|7/1=7
  reg ys97_o;  // 8:6|7/1=7
  reg ys98_o;  // 8:6|7/1=7
  reg ys99_o;  // 8:5|7/1=7
  reg ys100_o;  // 8:6|7/1=7
  reg ys101_o;  // 8:5|7/1=7
  reg ys102_o;  // 6:3|7/1=7
  reg ys103_o;  // 6:3|7/1=7
  reg ys104_o;  // 7:4|7/1=7
  reg ys105_o;  // 7:4|7/1=7
  reg ys106_o;  // 6:3|7/1=7
  reg ys107_o;  // 7:4|7/1=7
  reg ys108_o;  // 7:4|7/1=7
  reg ys109_o;  // 6:3|7/1=7
  reg ys110_o;  // 6:3|7/1=7
  reg ys111_o;  // 6:3|7/1=7
  reg ys112_o;  // 7:4|7/1=7
  reg ys113_o;  // 7:4|7/1=7
  reg ys114_o;  // 7:4|7/1=7
  reg ys115_o;  // 7:4|7/1=7
  reg ys116_o;  // 7:4|7/1=7
  reg ys117_o;  // 8:6|7/1=7
  reg ys118_o;  // 8:6|7/1=7
  reg ys119_o;  // 8:5|7/1=7
  reg ys120_o;  // 6:3|7/1=7
  reg ys121_o;  // 6:3|7/1=7
  reg ys122_o;  // 6:3|7/1=7
  reg ys123_o;  // 6:3|7/1=7
  reg ys124_o;  // 6:3|7/1=7
  reg ys125_o;  // 7:4|7/1=7
  reg ys126_o;  // 8:6|7/1=7
  reg ys127_o;  // 8:5|7/1=7
  reg ys128_o;  // 8:5|7/1=7
  reg ys129_o;  // 8:6|7/1=7
  reg ys130_o;  // 8:6|7/1=7
  reg ys131_o;  // 8:6|7/1=7
  reg ys132_o;  // 8:6|7/1=7
  reg ys133_o;  // 8:6|7/1=7
  reg ys134_o;  // 8:6|7/1=7
  reg ys135_o;  // 8:5|7/1=7
  reg ys136_o;  // 8:6|7/1=7
  reg ys137_o;  // 8:5|7/1=7
  reg ys138_o;  // 7:4|7/1=7
  reg ys139_o;  // 8:6|7/1=7
  reg ys140_o;  // 8:5|7/1=7
  reg ys141_o;  // 8:6|7/1=7
  reg ys142_o;  // 8:5|7/1=7
  reg ys143_o;  // 6:3|7/1=7
  reg ys144_o;  // 6:3|7/1=7
  reg ys145_o;  // 6:3|7/1=7
  reg ys146_o;  // 7:4|7/1=7
  reg ys147_o;  // 8:6|7/1=7
  reg ys148_o;  // 8:6|7/1=7
  reg ys149_o;  // 8:6|7/1=7
  reg ys150_o;  // 8:5|7/1=7
  reg ys151_o;  // 8:6|7/1=7
  reg ys152_o;  // 8:5|7/1=7
  reg ys153_o;  // 6:3|7/1=7
  reg ys154_o;  // 6:3|7/1=7
  reg ys155_o;  // 7:4|7/1=7
  reg ys156_o;  // 7:4|7/1=7
  reg ys157_o;  // 6:3|7/1=7
  reg ys158_o;  // 6:3|7/1=7
  reg ys159_o;  // 6:3|7/1=7
  reg ys160_o;  // 6:3|7/1=7
  reg ys161_o;  // 6:3|7/1=7
  reg ys162_o;  // 7:4|7/1=7
  reg ys163_o;  // 7:4|7/1=7
  reg ys164_o;  // 7:4|7/1=7
  reg ys165_o;  // 8:6|7/1=7
  reg ys166_o;  // 8:5|7/1=7
  reg ys167_o;  // 8:6|7/1=7
  reg ys168_o;  // 8:6|7/1=7
  reg ys169_o;  // 8:5|7/1=7
  reg ys170_o;  // 8:5|7/1=7
  reg ys171_o;  // 8:5|7/1=7
  reg ys172_o;  // 8:6|7/1=7
  reg ys173_o;  // 8:5|7/1=7
  reg ys174_o;  // 6:3|7/1=7
  reg ys175_o;  // 6:3|7/1=7
  reg ys176_o;  // 6:3|7/1=7
  reg ys177_o;  // 7:4|7/1=7
  reg ys178_o;  // 8:6|7/1=7
  reg ys179_o;  // 8:5|7/1=7
  reg ys180_o;  // 8:6|7/1=7
  reg ys181_o;  // 8:6|7/1=7
  reg ys182_o;  // 8:6|7/1=7
  reg ys183_o;  // 8:5|7/1=7

  wire ctre_cq0;
  wire ctre_cq1;
  wire ctre_cq2;
  wire ctre_cq3;
  wire ctre_cq4;
  wire ctre_cq5;
  wire ctre_cq6;
  wire ctre_cq7;
  wire ctre_cq8;
  wire ctre_cq9;
  wire ctre_cr0;
  wire ctre_cr1;
  wire ctre_cr2;
  wire ctre_cr3;
  wire ctre_cr4;
  wire ctre_cr5;
  wire ctre_cr6;
  wire ctre_cr7;
  wire ctre_cr8;
  wire ctre_cr9;
  wire ctre_dq;
  wire ctre_sq0;
  wire ctre_sq1;
  wire ctre_sq2;
  wire ctre_sq3;
  wire ctre_sq4;
  wire ctre_sq5;
  wire ctre_sq6;
  wire ctre_sq7;
  wire ctre_sq8;
  wire ctre_sq9;
  wire ctre_sr0;
  wire ctre_sr1;
  wire ctre_sr2;
  wire ctre_sr3;
  wire ctre_sr4;
  wire ctre_sr5;
  wire ctre_sr6;
  wire ctre_sr7;
  wire ctre_sr8;
  wire ctre_sr9;
  wire dn_o;
  wire jp;
  wire jpn;
  wire md;
  wire mdn;
  wire multm_compress_add3b_maj3b_or3b_wx0;
  wire multm_compress_add3b_maj3b_or3b_wx2;
  wire multm_compress_add3b_maj3b_or3b_wx3;
  wire multm_compress_add3b_maj3b_or3b_wx4;
  wire multm_compress_add3b_maj3b_or3b_wx5;
  wire multm_compress_add3b_maj3b_or3b_wx8;
  wire multm_compress_add3b_maj3b_or3b_wx9;
  wire multm_compress_add3b_maj3b_or3b_wx10;
  wire multm_compress_add3b_maj3b_or3b_wx11;
  wire multm_compress_add3b_maj3b_or3b_wx12;
  wire multm_compress_add3b_maj3b_or3b_wx13;
  wire multm_compress_add3b_maj3b_or3b_wx14;
  wire multm_compress_add3b_maj3b_or3b_wx15;
  wire multm_compress_add3b_maj3b_or3b_wx16;
  wire multm_compress_add3b_maj3b_or3b_wx17;
  wire multm_compress_add3b_maj3b_or3b_wx18;
  wire multm_compress_add3b_maj3b_or3b_wx19;
  wire multm_compress_add3b_maj3b_or3b_wx20;
  wire multm_compress_add3b_maj3b_or3b_wx21;
  wire multm_compress_add3b_maj3b_or3b_wx22;
  wire multm_compress_add3b_maj3b_or3b_wx23;
  wire multm_compress_add3b_maj3b_or3b_wx25;
  wire multm_compress_add3b_maj3b_or3b_wx26;
  wire multm_compress_add3b_maj3b_or3b_wx27;
  wire multm_compress_add3b_maj3b_or3b_wx28;
  wire multm_compress_add3b_maj3b_or3b_wx29;
  wire multm_compress_add3b_maj3b_or3b_wx30;
  wire multm_compress_add3b_maj3b_or3b_wx31;
  wire multm_compress_add3b_maj3b_or3b_wx32;
  wire multm_compress_add3b_maj3b_or3b_wx33;
  wire multm_compress_add3b_maj3b_or3b_wx34;
  wire multm_compress_add3b_maj3b_or3b_wx35;
  wire multm_compress_add3b_maj3b_or3b_wx36;
  wire multm_compress_add3b_maj3b_or3b_wx37;
  wire multm_compress_add3b_maj3b_or3b_wx38;
  wire multm_compress_add3b_maj3b_or3b_wx39;
  wire multm_compress_add3b_maj3b_or3b_wx40;
  wire multm_compress_add3b_maj3b_or3b_wx41;
  wire multm_compress_add3b_maj3b_or3b_wx44;
  wire multm_compress_add3b_maj3b_or3b_wx45;
  wire multm_compress_add3b_maj3b_or3b_wx46;
  wire multm_compress_add3b_maj3b_or3b_wx47;
  wire multm_compress_add3b_maj3b_or3b_wx48;
  wire multm_compress_add3b_maj3b_or3b_wx49;
  wire multm_compress_add3b_maj3b_or3b_wx50;
  wire multm_compress_add3b_maj3b_or3b_wx51;
  wire multm_compress_add3b_maj3b_or3b_wx52;
  wire multm_compress_add3b_maj3b_or3b_wx56;
  wire multm_compress_add3b_maj3b_or3b_wx57;
  wire multm_compress_add3b_maj3b_or3b_wx58;
  wire multm_compress_add3b_maj3b_or3b_wx59;
  wire multm_compress_add3b_maj3b_or3b_wx60;
  wire multm_compress_add3b_maj3b_or3b_wx61;
  wire multm_compress_add3b_maj3b_or3b_wx62;
  wire multm_compress_add3b_maj3b_or3b_wx63;
  wire multm_compress_add3b_maj3b_or3b_wx64;
  wire multm_compress_add3b_maj3b_or3b_wx65;
  wire multm_compress_add3b_maj3b_or3b_wx66;
  wire multm_compress_add3b_maj3b_or3b_wx67;
  wire multm_compress_add3b_maj3b_or3b_wx68;
  wire multm_compress_add3b_maj3b_or3b_wx69;
  wire multm_compress_add3b_maj3b_or3b_wx70;
  wire multm_compress_add3b_maj3b_or3b_wx71;
  wire multm_compress_add3b_maj3b_or3b_wx72;
  wire multm_compress_add3b_maj3b_or3b_wx73;
  wire multm_compress_add3b_maj3b_or3b_wx75;
  wire multm_compress_add3b_maj3b_or3b_wx76;
  wire multm_compress_add3b_maj3b_or3b_wx77;
  wire multm_compress_add3b_maj3b_or3b_wx78;
  wire multm_compress_add3b_maj3b_or3b_wx79;
  wire multm_compress_add3b_maj3b_or3b_wx80;
  wire multm_compress_add3b_maj3b_or3b_wx81;
  wire multm_compress_add3b_maj3b_or3b_wx82;
  wire multm_compress_add3b_maj3b_or3b_wx83;
  wire multm_compress_add3b_maj3b_or3b_wx84;
  wire multm_compress_add3b_maj3b_or3b_wx85;
  wire multm_compress_add3b_maj3b_or3b_wx86;
  wire multm_compress_add3b_maj3b_or3b_wx87;
  wire multm_compress_add3b_maj3b_or3b_wx88;
  wire multm_compress_add3b_maj3b_or3b_wx89;
  wire multm_compress_add3b_maj3b_or3b_wx90;
  wire multm_compress_add3b_maj3b_or3b_wx91;
  wire multm_compress_add3b_maj3b_or3b_wx92;
  wire multm_compress_add3b_maj3b_or3b_wx93;
  wire multm_compress_add3b_maj3b_or3b_wx94;
  wire multm_compress_add3b_maj3b_or3b_wx95;
  wire multm_compress_add3b_maj3b_or3b_wx96;
  wire multm_compress_add3b_maj3b_or3b_wx97;
  wire multm_compress_add3b_maj3b_or3b_wx98;
  wire multm_compress_add3b_maj3b_or3b_wx99;
  wire multm_compress_add3b_maj3b_or3b_wx100;
  wire multm_compress_add3b_maj3b_or3b_wx103;
  wire multm_compress_add3b_maj3b_or3b_wx104;
  wire multm_compress_add3b_maj3b_or3b_wx106;
  wire multm_compress_add3b_maj3b_or3b_wx107;
  wire multm_compress_add3b_maj3b_or3b_wx111;
  wire multm_compress_add3b_maj3b_or3b_wx112;
  wire multm_compress_add3b_maj3b_or3b_wx113;
  wire multm_compress_add3b_maj3b_or3b_wx114;
  wire multm_compress_add3b_maj3b_or3b_wx115;
  wire multm_compress_add3b_maj3b_or3b_wx116;
  wire multm_compress_add3b_maj3b_or3b_wx117;
  wire multm_compress_add3b_maj3b_or3b_wx118;
  wire multm_compress_add3b_maj3b_or3b_wx124;
  wire multm_compress_add3b_maj3b_or3b_wx125;
  wire multm_compress_add3b_maj3b_or3b_wx126;
  wire multm_compress_add3b_maj3b_or3b_wx127;
  wire multm_compress_add3b_maj3b_or3b_wx128;
  wire multm_compress_add3b_maj3b_or3b_wx129;
  wire multm_compress_add3b_maj3b_or3b_wx130;
  wire multm_compress_add3b_maj3b_or3b_wx131;
  wire multm_compress_add3b_maj3b_or3b_wx132;
  wire multm_compress_add3b_maj3b_or3b_wx133;
  wire multm_compress_add3b_maj3b_or3b_wx134;
  wire multm_compress_add3b_maj3b_or3b_wx135;
  wire multm_compress_add3b_maj3b_or3b_wx136;
  wire multm_compress_add3b_maj3b_or3b_wx137;
  wire multm_compress_add3b_maj3b_or3b_wx138;
  wire multm_compress_add3b_maj3b_or3b_wx139;
  wire multm_compress_add3b_maj3b_or3b_wx140;
  wire multm_compress_add3b_maj3b_or3b_wx141;
  wire multm_compress_add3b_maj3b_or3b_wx145;
  wire multm_compress_add3b_maj3b_or3b_wx146;
  wire multm_compress_add3b_maj3b_or3b_wx147;
  wire multm_compress_add3b_maj3b_or3b_wx148;
  wire multm_compress_add3b_maj3b_or3b_wx149;
  wire multm_compress_add3b_maj3b_or3b_wx150;
  wire multm_compress_add3b_maj3b_or3b_wx151;
  wire multm_compress_add3b_maj3b_or3b_wx154;
  wire multm_compress_add3b_maj3b_or3b_wx155;
  wire multm_compress_add3b_maj3b_or3b_wx161;
  wire multm_compress_add3b_maj3b_or3b_wx162;
  wire multm_compress_add3b_maj3b_or3b_wx163;
  wire multm_compress_add3b_maj3b_or3b_wx164;
  wire multm_compress_add3b_maj3b_or3b_wx165;
  wire multm_compress_add3b_maj3b_or3b_wx166;
  wire multm_compress_add3b_maj3b_or3b_wx167;
  wire multm_compress_add3b_maj3b_or3b_wx168;
  wire multm_compress_add3b_maj3b_or3b_wx169;
  wire multm_compress_add3b_maj3b_or3b_wx170;
  wire multm_compress_add3b_maj3b_or3b_wx171;
  wire multm_compress_add3b_maj3b_or3b_wx172;
  wire multm_compress_add3b_maj3b_or3b_wx176;
  wire multm_compress_add3b_maj3b_or3b_wx177;
  wire multm_compress_add3b_maj3b_or3b_wx178;
  wire multm_compress_add3b_maj3b_or3b_wx179;
  wire multm_compress_add3b_maj3b_or3b_wx180;
  wire multm_compress_add3b_maj3b_or3b_wx181;
  wire multm_compress_add3b_maj3b_or3b_wx182;
  wire multm_compress_add3b_maj3b_wx0;
  wire multm_compress_add3b_maj3b_wx2;
  wire multm_compress_add3b_maj3b_wx3;
  wire multm_compress_add3b_maj3b_wx4;
  wire multm_compress_add3b_maj3b_wx5;
  wire multm_compress_add3b_maj3b_wx8;
  wire multm_compress_add3b_maj3b_wx9;
  wire multm_compress_add3b_maj3b_wx10;
  wire multm_compress_add3b_maj3b_wx11;
  wire multm_compress_add3b_maj3b_wx12;
  wire multm_compress_add3b_maj3b_wx13;
  wire multm_compress_add3b_maj3b_wx14;
  wire multm_compress_add3b_maj3b_wx15;
  wire multm_compress_add3b_maj3b_wx16;
  wire multm_compress_add3b_maj3b_wx17;
  wire multm_compress_add3b_maj3b_wx18;
  wire multm_compress_add3b_maj3b_wx19;
  wire multm_compress_add3b_maj3b_wx20;
  wire multm_compress_add3b_maj3b_wx21;
  wire multm_compress_add3b_maj3b_wx22;
  wire multm_compress_add3b_maj3b_wx23;
  wire multm_compress_add3b_maj3b_wx25;
  wire multm_compress_add3b_maj3b_wx26;
  wire multm_compress_add3b_maj3b_wx27;
  wire multm_compress_add3b_maj3b_wx28;
  wire multm_compress_add3b_maj3b_wx29;
  wire multm_compress_add3b_maj3b_wx30;
  wire multm_compress_add3b_maj3b_wx31;
  wire multm_compress_add3b_maj3b_wx32;
  wire multm_compress_add3b_maj3b_wx33;
  wire multm_compress_add3b_maj3b_wx34;
  wire multm_compress_add3b_maj3b_wx35;
  wire multm_compress_add3b_maj3b_wx36;
  wire multm_compress_add3b_maj3b_wx37;
  wire multm_compress_add3b_maj3b_wx38;
  wire multm_compress_add3b_maj3b_wx39;
  wire multm_compress_add3b_maj3b_wx40;
  wire multm_compress_add3b_maj3b_wx41;
  wire multm_compress_add3b_maj3b_wx44;
  wire multm_compress_add3b_maj3b_wx45;
  wire multm_compress_add3b_maj3b_wx46;
  wire multm_compress_add3b_maj3b_wx47;
  wire multm_compress_add3b_maj3b_wx48;
  wire multm_compress_add3b_maj3b_wx49;
  wire multm_compress_add3b_maj3b_wx50;
  wire multm_compress_add3b_maj3b_wx51;
  wire multm_compress_add3b_maj3b_wx52;
  wire multm_compress_add3b_maj3b_wx56;
  wire multm_compress_add3b_maj3b_wx57;
  wire multm_compress_add3b_maj3b_wx58;
  wire multm_compress_add3b_maj3b_wx59;
  wire multm_compress_add3b_maj3b_wx60;
  wire multm_compress_add3b_maj3b_wx61;
  wire multm_compress_add3b_maj3b_wx62;
  wire multm_compress_add3b_maj3b_wx63;
  wire multm_compress_add3b_maj3b_wx64;
  wire multm_compress_add3b_maj3b_wx65;
  wire multm_compress_add3b_maj3b_wx66;
  wire multm_compress_add3b_maj3b_wx67;
  wire multm_compress_add3b_maj3b_wx68;
  wire multm_compress_add3b_maj3b_wx69;
  wire multm_compress_add3b_maj3b_wx70;
  wire multm_compress_add3b_maj3b_wx71;
  wire multm_compress_add3b_maj3b_wx72;
  wire multm_compress_add3b_maj3b_wx73;
  wire multm_compress_add3b_maj3b_wx75;
  wire multm_compress_add3b_maj3b_wx76;
  wire multm_compress_add3b_maj3b_wx77;
  wire multm_compress_add3b_maj3b_wx78;
  wire multm_compress_add3b_maj3b_wx79;
  wire multm_compress_add3b_maj3b_wx80;
  wire multm_compress_add3b_maj3b_wx81;
  wire multm_compress_add3b_maj3b_wx82;
  wire multm_compress_add3b_maj3b_wx83;
  wire multm_compress_add3b_maj3b_wx84;
  wire multm_compress_add3b_maj3b_wx85;
  wire multm_compress_add3b_maj3b_wx86;
  wire multm_compress_add3b_maj3b_wx87;
  wire multm_compress_add3b_maj3b_wx88;
  wire multm_compress_add3b_maj3b_wx89;
  wire multm_compress_add3b_maj3b_wx90;
  wire multm_compress_add3b_maj3b_wx91;
  wire multm_compress_add3b_maj3b_wx92;
  wire multm_compress_add3b_maj3b_wx93;
  wire multm_compress_add3b_maj3b_wx94;
  wire multm_compress_add3b_maj3b_wx95;
  wire multm_compress_add3b_maj3b_wx96;
  wire multm_compress_add3b_maj3b_wx97;
  wire multm_compress_add3b_maj3b_wx98;
  wire multm_compress_add3b_maj3b_wx99;
  wire multm_compress_add3b_maj3b_wx100;
  wire multm_compress_add3b_maj3b_wx103;
  wire multm_compress_add3b_maj3b_wx104;
  wire multm_compress_add3b_maj3b_wx106;
  wire multm_compress_add3b_maj3b_wx107;
  wire multm_compress_add3b_maj3b_wx111;
  wire multm_compress_add3b_maj3b_wx112;
  wire multm_compress_add3b_maj3b_wx113;
  wire multm_compress_add3b_maj3b_wx114;
  wire multm_compress_add3b_maj3b_wx115;
  wire multm_compress_add3b_maj3b_wx116;
  wire multm_compress_add3b_maj3b_wx117;
  wire multm_compress_add3b_maj3b_wx118;
  wire multm_compress_add3b_maj3b_wx124;
  wire multm_compress_add3b_maj3b_wx125;
  wire multm_compress_add3b_maj3b_wx126;
  wire multm_compress_add3b_maj3b_wx127;
  wire multm_compress_add3b_maj3b_wx128;
  wire multm_compress_add3b_maj3b_wx129;
  wire multm_compress_add3b_maj3b_wx130;
  wire multm_compress_add3b_maj3b_wx131;
  wire multm_compress_add3b_maj3b_wx132;
  wire multm_compress_add3b_maj3b_wx133;
  wire multm_compress_add3b_maj3b_wx134;
  wire multm_compress_add3b_maj3b_wx135;
  wire multm_compress_add3b_maj3b_wx136;
  wire multm_compress_add3b_maj3b_wx137;
  wire multm_compress_add3b_maj3b_wx138;
  wire multm_compress_add3b_maj3b_wx139;
  wire multm_compress_add3b_maj3b_wx140;
  wire multm_compress_add3b_maj3b_wx141;
  wire multm_compress_add3b_maj3b_wx145;
  wire multm_compress_add3b_maj3b_wx146;
  wire multm_compress_add3b_maj3b_wx147;
  wire multm_compress_add3b_maj3b_wx148;
  wire multm_compress_add3b_maj3b_wx149;
  wire multm_compress_add3b_maj3b_wx150;
  wire multm_compress_add3b_maj3b_wx151;
  wire multm_compress_add3b_maj3b_wx154;
  wire multm_compress_add3b_maj3b_wx155;
  wire multm_compress_add3b_maj3b_wx161;
  wire multm_compress_add3b_maj3b_wx162;
  wire multm_compress_add3b_maj3b_wx163;
  wire multm_compress_add3b_maj3b_wx164;
  wire multm_compress_add3b_maj3b_wx165;
  wire multm_compress_add3b_maj3b_wx166;
  wire multm_compress_add3b_maj3b_wx167;
  wire multm_compress_add3b_maj3b_wx168;
  wire multm_compress_add3b_maj3b_wx169;
  wire multm_compress_add3b_maj3b_wx170;
  wire multm_compress_add3b_maj3b_wx171;
  wire multm_compress_add3b_maj3b_wx172;
  wire multm_compress_add3b_maj3b_wx176;
  wire multm_compress_add3b_maj3b_wx177;
  wire multm_compress_add3b_maj3b_wx178;
  wire multm_compress_add3b_maj3b_wx179;
  wire multm_compress_add3b_maj3b_wx180;
  wire multm_compress_add3b_maj3b_wx181;
  wire multm_compress_add3b_maj3b_wx182;
  wire multm_compress_add3b_maj3b_wy0;
  wire multm_compress_add3b_maj3b_wy2;
  wire multm_compress_add3b_maj3b_wy3;
  wire multm_compress_add3b_maj3b_wy4;
  wire multm_compress_add3b_maj3b_wy5;
  wire multm_compress_add3b_maj3b_wy8;
  wire multm_compress_add3b_maj3b_wy9;
  wire multm_compress_add3b_maj3b_wy10;
  wire multm_compress_add3b_maj3b_wy11;
  wire multm_compress_add3b_maj3b_wy12;
  wire multm_compress_add3b_maj3b_wy13;
  wire multm_compress_add3b_maj3b_wy14;
  wire multm_compress_add3b_maj3b_wy15;
  wire multm_compress_add3b_maj3b_wy16;
  wire multm_compress_add3b_maj3b_wy17;
  wire multm_compress_add3b_maj3b_wy18;
  wire multm_compress_add3b_maj3b_wy19;
  wire multm_compress_add3b_maj3b_wy20;
  wire multm_compress_add3b_maj3b_wy21;
  wire multm_compress_add3b_maj3b_wy22;
  wire multm_compress_add3b_maj3b_wy23;
  wire multm_compress_add3b_maj3b_wy25;
  wire multm_compress_add3b_maj3b_wy26;
  wire multm_compress_add3b_maj3b_wy27;
  wire multm_compress_add3b_maj3b_wy28;
  wire multm_compress_add3b_maj3b_wy29;
  wire multm_compress_add3b_maj3b_wy30;
  wire multm_compress_add3b_maj3b_wy31;
  wire multm_compress_add3b_maj3b_wy32;
  wire multm_compress_add3b_maj3b_wy33;
  wire multm_compress_add3b_maj3b_wy34;
  wire multm_compress_add3b_maj3b_wy35;
  wire multm_compress_add3b_maj3b_wy36;
  wire multm_compress_add3b_maj3b_wy37;
  wire multm_compress_add3b_maj3b_wy38;
  wire multm_compress_add3b_maj3b_wy39;
  wire multm_compress_add3b_maj3b_wy40;
  wire multm_compress_add3b_maj3b_wy41;
  wire multm_compress_add3b_maj3b_wy44;
  wire multm_compress_add3b_maj3b_wy45;
  wire multm_compress_add3b_maj3b_wy46;
  wire multm_compress_add3b_maj3b_wy47;
  wire multm_compress_add3b_maj3b_wy48;
  wire multm_compress_add3b_maj3b_wy49;
  wire multm_compress_add3b_maj3b_wy50;
  wire multm_compress_add3b_maj3b_wy51;
  wire multm_compress_add3b_maj3b_wy52;
  wire multm_compress_add3b_maj3b_wy56;
  wire multm_compress_add3b_maj3b_wy57;
  wire multm_compress_add3b_maj3b_wy58;
  wire multm_compress_add3b_maj3b_wy59;
  wire multm_compress_add3b_maj3b_wy60;
  wire multm_compress_add3b_maj3b_wy61;
  wire multm_compress_add3b_maj3b_wy62;
  wire multm_compress_add3b_maj3b_wy63;
  wire multm_compress_add3b_maj3b_wy64;
  wire multm_compress_add3b_maj3b_wy65;
  wire multm_compress_add3b_maj3b_wy66;
  wire multm_compress_add3b_maj3b_wy67;
  wire multm_compress_add3b_maj3b_wy68;
  wire multm_compress_add3b_maj3b_wy69;
  wire multm_compress_add3b_maj3b_wy70;
  wire multm_compress_add3b_maj3b_wy71;
  wire multm_compress_add3b_maj3b_wy72;
  wire multm_compress_add3b_maj3b_wy73;
  wire multm_compress_add3b_maj3b_wy75;
  wire multm_compress_add3b_maj3b_wy76;
  wire multm_compress_add3b_maj3b_wy77;
  wire multm_compress_add3b_maj3b_wy78;
  wire multm_compress_add3b_maj3b_wy79;
  wire multm_compress_add3b_maj3b_wy80;
  wire multm_compress_add3b_maj3b_wy81;
  wire multm_compress_add3b_maj3b_wy82;
  wire multm_compress_add3b_maj3b_wy83;
  wire multm_compress_add3b_maj3b_wy84;
  wire multm_compress_add3b_maj3b_wy85;
  wire multm_compress_add3b_maj3b_wy86;
  wire multm_compress_add3b_maj3b_wy87;
  wire multm_compress_add3b_maj3b_wy88;
  wire multm_compress_add3b_maj3b_wy89;
  wire multm_compress_add3b_maj3b_wy90;
  wire multm_compress_add3b_maj3b_wy91;
  wire multm_compress_add3b_maj3b_wy92;
  wire multm_compress_add3b_maj3b_wy93;
  wire multm_compress_add3b_maj3b_wy94;
  wire multm_compress_add3b_maj3b_wy95;
  wire multm_compress_add3b_maj3b_wy96;
  wire multm_compress_add3b_maj3b_wy97;
  wire multm_compress_add3b_maj3b_wy98;
  wire multm_compress_add3b_maj3b_wy99;
  wire multm_compress_add3b_maj3b_wy100;
  wire multm_compress_add3b_maj3b_wy103;
  wire multm_compress_add3b_maj3b_wy104;
  wire multm_compress_add3b_maj3b_wy106;
  wire multm_compress_add3b_maj3b_wy107;
  wire multm_compress_add3b_maj3b_wy111;
  wire multm_compress_add3b_maj3b_wy112;
  wire multm_compress_add3b_maj3b_wy113;
  wire multm_compress_add3b_maj3b_wy114;
  wire multm_compress_add3b_maj3b_wy115;
  wire multm_compress_add3b_maj3b_wy116;
  wire multm_compress_add3b_maj3b_wy117;
  wire multm_compress_add3b_maj3b_wy118;
  wire multm_compress_add3b_maj3b_wy124;
  wire multm_compress_add3b_maj3b_wy125;
  wire multm_compress_add3b_maj3b_wy126;
  wire multm_compress_add3b_maj3b_wy127;
  wire multm_compress_add3b_maj3b_wy128;
  wire multm_compress_add3b_maj3b_wy129;
  wire multm_compress_add3b_maj3b_wy130;
  wire multm_compress_add3b_maj3b_wy131;
  wire multm_compress_add3b_maj3b_wy132;
  wire multm_compress_add3b_maj3b_wy133;
  wire multm_compress_add3b_maj3b_wy134;
  wire multm_compress_add3b_maj3b_wy135;
  wire multm_compress_add3b_maj3b_wy136;
  wire multm_compress_add3b_maj3b_wy137;
  wire multm_compress_add3b_maj3b_wy138;
  wire multm_compress_add3b_maj3b_wy139;
  wire multm_compress_add3b_maj3b_wy140;
  wire multm_compress_add3b_maj3b_wy141;
  wire multm_compress_add3b_maj3b_wy145;
  wire multm_compress_add3b_maj3b_wy146;
  wire multm_compress_add3b_maj3b_wy147;
  wire multm_compress_add3b_maj3b_wy148;
  wire multm_compress_add3b_maj3b_wy149;
  wire multm_compress_add3b_maj3b_wy150;
  wire multm_compress_add3b_maj3b_wy151;
  wire multm_compress_add3b_maj3b_wy154;
  wire multm_compress_add3b_maj3b_wy155;
  wire multm_compress_add3b_maj3b_wy161;
  wire multm_compress_add3b_maj3b_wy162;
  wire multm_compress_add3b_maj3b_wy163;
  wire multm_compress_add3b_maj3b_wy164;
  wire multm_compress_add3b_maj3b_wy165;
  wire multm_compress_add3b_maj3b_wy166;
  wire multm_compress_add3b_maj3b_wy167;
  wire multm_compress_add3b_maj3b_wy168;
  wire multm_compress_add3b_maj3b_wy169;
  wire multm_compress_add3b_maj3b_wy170;
  wire multm_compress_add3b_maj3b_wy171;
  wire multm_compress_add3b_maj3b_wy172;
  wire multm_compress_add3b_maj3b_wy176;
  wire multm_compress_add3b_maj3b_wy177;
  wire multm_compress_add3b_maj3b_wy178;
  wire multm_compress_add3b_maj3b_wy179;
  wire multm_compress_add3b_maj3b_wy180;
  wire multm_compress_add3b_maj3b_wy181;
  wire multm_compress_add3b_maj3b_wy182;
  wire multm_compress_add3b_maj3b_xy0;
  wire multm_compress_add3b_maj3b_xy2;
  wire multm_compress_add3b_maj3b_xy3;
  wire multm_compress_add3b_maj3b_xy4;
  wire multm_compress_add3b_maj3b_xy5;
  wire multm_compress_add3b_maj3b_xy8;
  wire multm_compress_add3b_maj3b_xy9;
  wire multm_compress_add3b_maj3b_xy10;
  wire multm_compress_add3b_maj3b_xy11;
  wire multm_compress_add3b_maj3b_xy12;
  wire multm_compress_add3b_maj3b_xy13;
  wire multm_compress_add3b_maj3b_xy14;
  wire multm_compress_add3b_maj3b_xy15;
  wire multm_compress_add3b_maj3b_xy16;
  wire multm_compress_add3b_maj3b_xy17;
  wire multm_compress_add3b_maj3b_xy18;
  wire multm_compress_add3b_maj3b_xy19;
  wire multm_compress_add3b_maj3b_xy20;
  wire multm_compress_add3b_maj3b_xy21;
  wire multm_compress_add3b_maj3b_xy22;
  wire multm_compress_add3b_maj3b_xy23;
  wire multm_compress_add3b_maj3b_xy25;
  wire multm_compress_add3b_maj3b_xy26;
  wire multm_compress_add3b_maj3b_xy27;
  wire multm_compress_add3b_maj3b_xy28;
  wire multm_compress_add3b_maj3b_xy29;
  wire multm_compress_add3b_maj3b_xy30;
  wire multm_compress_add3b_maj3b_xy31;
  wire multm_compress_add3b_maj3b_xy32;
  wire multm_compress_add3b_maj3b_xy33;
  wire multm_compress_add3b_maj3b_xy34;
  wire multm_compress_add3b_maj3b_xy35;
  wire multm_compress_add3b_maj3b_xy36;
  wire multm_compress_add3b_maj3b_xy37;
  wire multm_compress_add3b_maj3b_xy38;
  wire multm_compress_add3b_maj3b_xy39;
  wire multm_compress_add3b_maj3b_xy40;
  wire multm_compress_add3b_maj3b_xy41;
  wire multm_compress_add3b_maj3b_xy44;
  wire multm_compress_add3b_maj3b_xy45;
  wire multm_compress_add3b_maj3b_xy46;
  wire multm_compress_add3b_maj3b_xy47;
  wire multm_compress_add3b_maj3b_xy48;
  wire multm_compress_add3b_maj3b_xy49;
  wire multm_compress_add3b_maj3b_xy50;
  wire multm_compress_add3b_maj3b_xy51;
  wire multm_compress_add3b_maj3b_xy52;
  wire multm_compress_add3b_maj3b_xy56;
  wire multm_compress_add3b_maj3b_xy57;
  wire multm_compress_add3b_maj3b_xy58;
  wire multm_compress_add3b_maj3b_xy59;
  wire multm_compress_add3b_maj3b_xy60;
  wire multm_compress_add3b_maj3b_xy61;
  wire multm_compress_add3b_maj3b_xy62;
  wire multm_compress_add3b_maj3b_xy63;
  wire multm_compress_add3b_maj3b_xy64;
  wire multm_compress_add3b_maj3b_xy65;
  wire multm_compress_add3b_maj3b_xy66;
  wire multm_compress_add3b_maj3b_xy67;
  wire multm_compress_add3b_maj3b_xy68;
  wire multm_compress_add3b_maj3b_xy69;
  wire multm_compress_add3b_maj3b_xy70;
  wire multm_compress_add3b_maj3b_xy71;
  wire multm_compress_add3b_maj3b_xy72;
  wire multm_compress_add3b_maj3b_xy73;
  wire multm_compress_add3b_maj3b_xy75;
  wire multm_compress_add3b_maj3b_xy76;
  wire multm_compress_add3b_maj3b_xy77;
  wire multm_compress_add3b_maj3b_xy78;
  wire multm_compress_add3b_maj3b_xy79;
  wire multm_compress_add3b_maj3b_xy80;
  wire multm_compress_add3b_maj3b_xy81;
  wire multm_compress_add3b_maj3b_xy82;
  wire multm_compress_add3b_maj3b_xy83;
  wire multm_compress_add3b_maj3b_xy84;
  wire multm_compress_add3b_maj3b_xy85;
  wire multm_compress_add3b_maj3b_xy86;
  wire multm_compress_add3b_maj3b_xy87;
  wire multm_compress_add3b_maj3b_xy88;
  wire multm_compress_add3b_maj3b_xy89;
  wire multm_compress_add3b_maj3b_xy90;
  wire multm_compress_add3b_maj3b_xy91;
  wire multm_compress_add3b_maj3b_xy92;
  wire multm_compress_add3b_maj3b_xy93;
  wire multm_compress_add3b_maj3b_xy94;
  wire multm_compress_add3b_maj3b_xy95;
  wire multm_compress_add3b_maj3b_xy96;
  wire multm_compress_add3b_maj3b_xy97;
  wire multm_compress_add3b_maj3b_xy98;
  wire multm_compress_add3b_maj3b_xy99;
  wire multm_compress_add3b_maj3b_xy100;
  wire multm_compress_add3b_maj3b_xy103;
  wire multm_compress_add3b_maj3b_xy104;
  wire multm_compress_add3b_maj3b_xy106;
  wire multm_compress_add3b_maj3b_xy107;
  wire multm_compress_add3b_maj3b_xy111;
  wire multm_compress_add3b_maj3b_xy112;
  wire multm_compress_add3b_maj3b_xy113;
  wire multm_compress_add3b_maj3b_xy114;
  wire multm_compress_add3b_maj3b_xy115;
  wire multm_compress_add3b_maj3b_xy116;
  wire multm_compress_add3b_maj3b_xy117;
  wire multm_compress_add3b_maj3b_xy118;
  wire multm_compress_add3b_maj3b_xy124;
  wire multm_compress_add3b_maj3b_xy125;
  wire multm_compress_add3b_maj3b_xy126;
  wire multm_compress_add3b_maj3b_xy127;
  wire multm_compress_add3b_maj3b_xy128;
  wire multm_compress_add3b_maj3b_xy129;
  wire multm_compress_add3b_maj3b_xy130;
  wire multm_compress_add3b_maj3b_xy131;
  wire multm_compress_add3b_maj3b_xy132;
  wire multm_compress_add3b_maj3b_xy133;
  wire multm_compress_add3b_maj3b_xy134;
  wire multm_compress_add3b_maj3b_xy135;
  wire multm_compress_add3b_maj3b_xy136;
  wire multm_compress_add3b_maj3b_xy137;
  wire multm_compress_add3b_maj3b_xy138;
  wire multm_compress_add3b_maj3b_xy139;
  wire multm_compress_add3b_maj3b_xy140;
  wire multm_compress_add3b_maj3b_xy141;
  wire multm_compress_add3b_maj3b_xy145;
  wire multm_compress_add3b_maj3b_xy146;
  wire multm_compress_add3b_maj3b_xy147;
  wire multm_compress_add3b_maj3b_xy148;
  wire multm_compress_add3b_maj3b_xy149;
  wire multm_compress_add3b_maj3b_xy150;
  wire multm_compress_add3b_maj3b_xy151;
  wire multm_compress_add3b_maj3b_xy154;
  wire multm_compress_add3b_maj3b_xy155;
  wire multm_compress_add3b_maj3b_xy161;
  wire multm_compress_add3b_maj3b_xy162;
  wire multm_compress_add3b_maj3b_xy163;
  wire multm_compress_add3b_maj3b_xy164;
  wire multm_compress_add3b_maj3b_xy165;
  wire multm_compress_add3b_maj3b_xy166;
  wire multm_compress_add3b_maj3b_xy167;
  wire multm_compress_add3b_maj3b_xy168;
  wire multm_compress_add3b_maj3b_xy169;
  wire multm_compress_add3b_maj3b_xy170;
  wire multm_compress_add3b_maj3b_xy171;
  wire multm_compress_add3b_maj3b_xy172;
  wire multm_compress_add3b_maj3b_xy176;
  wire multm_compress_add3b_maj3b_xy177;
  wire multm_compress_add3b_maj3b_xy178;
  wire multm_compress_add3b_maj3b_xy179;
  wire multm_compress_add3b_maj3b_xy180;
  wire multm_compress_add3b_maj3b_xy181;
  wire multm_compress_add3b_maj3b_xy182;
  wire multm_compress_add3b_xor3b_wx0;
  wire multm_compress_add3b_xor3b_wx2;
  wire multm_compress_add3b_xor3b_wx3;
  wire multm_compress_add3b_xor3b_wx4;
  wire multm_compress_add3b_xor3b_wx5;
  wire multm_compress_add3b_xor3b_wx8;
  wire multm_compress_add3b_xor3b_wx9;
  wire multm_compress_add3b_xor3b_wx10;
  wire multm_compress_add3b_xor3b_wx11;
  wire multm_compress_add3b_xor3b_wx12;
  wire multm_compress_add3b_xor3b_wx13;
  wire multm_compress_add3b_xor3b_wx14;
  wire multm_compress_add3b_xor3b_wx15;
  wire multm_compress_add3b_xor3b_wx16;
  wire multm_compress_add3b_xor3b_wx17;
  wire multm_compress_add3b_xor3b_wx18;
  wire multm_compress_add3b_xor3b_wx19;
  wire multm_compress_add3b_xor3b_wx20;
  wire multm_compress_add3b_xor3b_wx21;
  wire multm_compress_add3b_xor3b_wx22;
  wire multm_compress_add3b_xor3b_wx23;
  wire multm_compress_add3b_xor3b_wx25;
  wire multm_compress_add3b_xor3b_wx26;
  wire multm_compress_add3b_xor3b_wx27;
  wire multm_compress_add3b_xor3b_wx28;
  wire multm_compress_add3b_xor3b_wx29;
  wire multm_compress_add3b_xor3b_wx30;
  wire multm_compress_add3b_xor3b_wx31;
  wire multm_compress_add3b_xor3b_wx32;
  wire multm_compress_add3b_xor3b_wx33;
  wire multm_compress_add3b_xor3b_wx34;
  wire multm_compress_add3b_xor3b_wx35;
  wire multm_compress_add3b_xor3b_wx36;
  wire multm_compress_add3b_xor3b_wx37;
  wire multm_compress_add3b_xor3b_wx38;
  wire multm_compress_add3b_xor3b_wx39;
  wire multm_compress_add3b_xor3b_wx40;
  wire multm_compress_add3b_xor3b_wx41;
  wire multm_compress_add3b_xor3b_wx44;
  wire multm_compress_add3b_xor3b_wx45;
  wire multm_compress_add3b_xor3b_wx46;
  wire multm_compress_add3b_xor3b_wx47;
  wire multm_compress_add3b_xor3b_wx48;
  wire multm_compress_add3b_xor3b_wx49;
  wire multm_compress_add3b_xor3b_wx50;
  wire multm_compress_add3b_xor3b_wx51;
  wire multm_compress_add3b_xor3b_wx52;
  wire multm_compress_add3b_xor3b_wx56;
  wire multm_compress_add3b_xor3b_wx57;
  wire multm_compress_add3b_xor3b_wx58;
  wire multm_compress_add3b_xor3b_wx59;
  wire multm_compress_add3b_xor3b_wx60;
  wire multm_compress_add3b_xor3b_wx61;
  wire multm_compress_add3b_xor3b_wx62;
  wire multm_compress_add3b_xor3b_wx63;
  wire multm_compress_add3b_xor3b_wx64;
  wire multm_compress_add3b_xor3b_wx65;
  wire multm_compress_add3b_xor3b_wx66;
  wire multm_compress_add3b_xor3b_wx67;
  wire multm_compress_add3b_xor3b_wx68;
  wire multm_compress_add3b_xor3b_wx69;
  wire multm_compress_add3b_xor3b_wx70;
  wire multm_compress_add3b_xor3b_wx71;
  wire multm_compress_add3b_xor3b_wx72;
  wire multm_compress_add3b_xor3b_wx73;
  wire multm_compress_add3b_xor3b_wx75;
  wire multm_compress_add3b_xor3b_wx76;
  wire multm_compress_add3b_xor3b_wx77;
  wire multm_compress_add3b_xor3b_wx78;
  wire multm_compress_add3b_xor3b_wx79;
  wire multm_compress_add3b_xor3b_wx80;
  wire multm_compress_add3b_xor3b_wx81;
  wire multm_compress_add3b_xor3b_wx82;
  wire multm_compress_add3b_xor3b_wx83;
  wire multm_compress_add3b_xor3b_wx84;
  wire multm_compress_add3b_xor3b_wx85;
  wire multm_compress_add3b_xor3b_wx86;
  wire multm_compress_add3b_xor3b_wx87;
  wire multm_compress_add3b_xor3b_wx88;
  wire multm_compress_add3b_xor3b_wx89;
  wire multm_compress_add3b_xor3b_wx90;
  wire multm_compress_add3b_xor3b_wx91;
  wire multm_compress_add3b_xor3b_wx92;
  wire multm_compress_add3b_xor3b_wx93;
  wire multm_compress_add3b_xor3b_wx94;
  wire multm_compress_add3b_xor3b_wx95;
  wire multm_compress_add3b_xor3b_wx96;
  wire multm_compress_add3b_xor3b_wx97;
  wire multm_compress_add3b_xor3b_wx98;
  wire multm_compress_add3b_xor3b_wx99;
  wire multm_compress_add3b_xor3b_wx100;
  wire multm_compress_add3b_xor3b_wx103;
  wire multm_compress_add3b_xor3b_wx104;
  wire multm_compress_add3b_xor3b_wx106;
  wire multm_compress_add3b_xor3b_wx107;
  wire multm_compress_add3b_xor3b_wx111;
  wire multm_compress_add3b_xor3b_wx112;
  wire multm_compress_add3b_xor3b_wx113;
  wire multm_compress_add3b_xor3b_wx114;
  wire multm_compress_add3b_xor3b_wx115;
  wire multm_compress_add3b_xor3b_wx116;
  wire multm_compress_add3b_xor3b_wx117;
  wire multm_compress_add3b_xor3b_wx118;
  wire multm_compress_add3b_xor3b_wx124;
  wire multm_compress_add3b_xor3b_wx125;
  wire multm_compress_add3b_xor3b_wx126;
  wire multm_compress_add3b_xor3b_wx127;
  wire multm_compress_add3b_xor3b_wx128;
  wire multm_compress_add3b_xor3b_wx129;
  wire multm_compress_add3b_xor3b_wx130;
  wire multm_compress_add3b_xor3b_wx131;
  wire multm_compress_add3b_xor3b_wx132;
  wire multm_compress_add3b_xor3b_wx133;
  wire multm_compress_add3b_xor3b_wx134;
  wire multm_compress_add3b_xor3b_wx135;
  wire multm_compress_add3b_xor3b_wx136;
  wire multm_compress_add3b_xor3b_wx137;
  wire multm_compress_add3b_xor3b_wx138;
  wire multm_compress_add3b_xor3b_wx139;
  wire multm_compress_add3b_xor3b_wx140;
  wire multm_compress_add3b_xor3b_wx141;
  wire multm_compress_add3b_xor3b_wx145;
  wire multm_compress_add3b_xor3b_wx146;
  wire multm_compress_add3b_xor3b_wx147;
  wire multm_compress_add3b_xor3b_wx148;
  wire multm_compress_add3b_xor3b_wx149;
  wire multm_compress_add3b_xor3b_wx150;
  wire multm_compress_add3b_xor3b_wx151;
  wire multm_compress_add3b_xor3b_wx154;
  wire multm_compress_add3b_xor3b_wx155;
  wire multm_compress_add3b_xor3b_wx161;
  wire multm_compress_add3b_xor3b_wx162;
  wire multm_compress_add3b_xor3b_wx163;
  wire multm_compress_add3b_xor3b_wx164;
  wire multm_compress_add3b_xor3b_wx165;
  wire multm_compress_add3b_xor3b_wx166;
  wire multm_compress_add3b_xor3b_wx167;
  wire multm_compress_add3b_xor3b_wx168;
  wire multm_compress_add3b_xor3b_wx169;
  wire multm_compress_add3b_xor3b_wx170;
  wire multm_compress_add3b_xor3b_wx171;
  wire multm_compress_add3b_xor3b_wx172;
  wire multm_compress_add3b_xor3b_wx176;
  wire multm_compress_add3b_xor3b_wx177;
  wire multm_compress_add3b_xor3b_wx178;
  wire multm_compress_add3b_xor3b_wx179;
  wire multm_compress_add3b_xor3b_wx180;
  wire multm_compress_add3b_xor3b_wx181;
  wire multm_compress_add3b_xor3b_wx182;
  wire multm_compress_nc;
  wire multm_compress_nct;
  wire multm_compress_ns;
  wire multm_compress_rn4;
  wire multm_compress_rn5;
  wire multm_compress_rn6;
  wire multm_compress_rn15;
  wire multm_compress_rn20;
  wire multm_compress_rnh4;
  wire multm_ctrp_ctr_cq0;
  wire multm_ctrp_ctr_cq1;
  wire multm_ctrp_ctr_cq2;
  wire multm_ctrp_ctr_cq3;
  wire multm_ctrp_ctr_cq4;
  wire multm_ctrp_ctr_cq5;
  wire multm_ctrp_ctr_cq6;
  wire multm_ctrp_ctr_cq7;
  wire multm_ctrp_ctr_cr0;
  wire multm_ctrp_ctr_cr1;
  wire multm_ctrp_ctr_cr2;
  wire multm_ctrp_ctr_cr3;
  wire multm_ctrp_ctr_cr4;
  wire multm_ctrp_ctr_cr5;
  wire multm_ctrp_ctr_cr6;
  wire multm_ctrp_ctr_cr7;
  wire multm_ctrp_ctr_dq;
  wire multm_ctrp_ctr_sq0;
  wire multm_ctrp_ctr_sq1;
  wire multm_ctrp_ctr_sq2;
  wire multm_ctrp_ctr_sq3;
  wire multm_ctrp_ctr_sq4;
  wire multm_ctrp_ctr_sq5;
  wire multm_ctrp_ctr_sq6;
  wire multm_ctrp_ctr_sr0;
  wire multm_ctrp_ctr_sr1;
  wire multm_ctrp_ctr_sr2;
  wire multm_ctrp_ctr_sr3;
  wire multm_ctrp_ctr_sr4;
  wire multm_ctrp_ctr_sr5;
  wire multm_ctrp_ctr_sr6;
  wire multm_ctrp_ds;
  wire multm_ctrp_pulse_xn;
  wire multm_pc0;
  wire multm_pc1;
  wire multm_pc2;
  wire multm_pc3;
  wire multm_pc4;
  wire multm_pc5;
  wire multm_pc6;
  wire multm_pc7;
  wire multm_pc8;
  wire multm_pc9;
  wire multm_pc11;
  wire multm_pc12;
  wire multm_pc13;
  wire multm_pc14;
  wire multm_pc15;
  wire multm_pc16;
  wire multm_pc17;
  wire multm_pc18;
  wire multm_pc19;
  wire multm_pc20;
  wire multm_pc21;
  wire multm_pc22;
  wire multm_pc23;
  wire multm_pc24;
  wire multm_pc25;
  wire multm_pc26;
  wire multm_pc27;
  wire multm_pc28;
  wire multm_pc29;
  wire multm_pc30;
  wire multm_pc31;
  wire multm_pc32;
  wire multm_pc33;
  wire multm_pc34;
  wire multm_pc35;
  wire multm_pc36;
  wire multm_pc37;
  wire multm_pc38;
  wire multm_pc39;
  wire multm_pc40;
  wire multm_pc41;
  wire multm_pc42;
  wire multm_pc43;
  wire multm_pc44;
  wire multm_pc45;
  wire multm_pc46;
  wire multm_pc47;
  wire multm_pc48;
  wire multm_pc49;
  wire multm_pc50;
  wire multm_pc51;
  wire multm_pc52;
  wire multm_pc53;
  wire multm_pc54;
  wire multm_pc55;
  wire multm_pc56;
  wire multm_pc57;
  wire multm_pc58;
  wire multm_pc59;
  wire multm_pc60;
  wire multm_pc61;
  wire multm_pc62;
  wire multm_pc63;
  wire multm_pc64;
  wire multm_pc65;
  wire multm_pc66;
  wire multm_pc67;
  wire multm_pc68;
  wire multm_pc69;
  wire multm_pc70;
  wire multm_pc71;
  wire multm_pc72;
  wire multm_pc73;
  wire multm_pc74;
  wire multm_pc75;
  wire multm_pc76;
  wire multm_pc77;
  wire multm_pc78;
  wire multm_pc79;
  wire multm_pc80;
  wire multm_pc81;
  wire multm_pc82;
  wire multm_pc83;
  wire multm_pc84;
  wire multm_pc85;
  wire multm_pc86;
  wire multm_pc87;
  wire multm_pc88;
  wire multm_pc89;
  wire multm_pc90;
  wire multm_pc91;
  wire multm_pc92;
  wire multm_pc93;
  wire multm_pc94;
  wire multm_pc95;
  wire multm_pc96;
  wire multm_pc97;
  wire multm_pc98;
  wire multm_pc99;
  wire multm_pc100;
  wire multm_pc101;
  wire multm_pc102;
  wire multm_pc103;
  wire multm_pc104;
  wire multm_pc105;
  wire multm_pc106;
  wire multm_pc107;
  wire multm_pc108;
  wire multm_pc109;
  wire multm_pc110;
  wire multm_pc111;
  wire multm_pc112;
  wire multm_pc113;
  wire multm_pc114;
  wire multm_pc115;
  wire multm_pc116;
  wire multm_pc117;
  wire multm_pc118;
  wire multm_pc119;
  wire multm_pc120;
  wire multm_pc121;
  wire multm_pc122;
  wire multm_pc123;
  wire multm_pc124;
  wire multm_pc125;
  wire multm_pc126;
  wire multm_pc127;
  wire multm_pc128;
  wire multm_pc129;
  wire multm_pc130;
  wire multm_pc131;
  wire multm_pc132;
  wire multm_pc133;
  wire multm_pc134;
  wire multm_pc135;
  wire multm_pc136;
  wire multm_pc137;
  wire multm_pc138;
  wire multm_pc139;
  wire multm_pc140;
  wire multm_pc141;
  wire multm_pc142;
  wire multm_pc143;
  wire multm_pc144;
  wire multm_pc145;
  wire multm_pc146;
  wire multm_pc147;
  wire multm_pc148;
  wire multm_pc149;
  wire multm_pc150;
  wire multm_pc151;
  wire multm_pc152;
  wire multm_pc153;
  wire multm_pc154;
  wire multm_pc155;
  wire multm_pc156;
  wire multm_pc157;
  wire multm_pc158;
  wire multm_pc159;
  wire multm_pc160;
  wire multm_pc161;
  wire multm_pc162;
  wire multm_pc163;
  wire multm_pc164;
  wire multm_pc165;
  wire multm_pc166;
  wire multm_pc167;
  wire multm_pc168;
  wire multm_pc169;
  wire multm_pc170;
  wire multm_pc171;
  wire multm_pc172;
  wire multm_pc173;
  wire multm_pc174;
  wire multm_pc175;
  wire multm_pc176;
  wire multm_pc177;
  wire multm_pc178;
  wire multm_pc179;
  wire multm_pc180;
  wire multm_pc181;
  wire multm_pc182;
  wire multm_pc183;
  wire multm_pc184;
  wire multm_ps0;
  wire multm_ps1;
  wire multm_ps2;
  wire multm_ps3;
  wire multm_ps4;
  wire multm_ps5;
  wire multm_ps6;
  wire multm_ps7;
  wire multm_ps8;
  wire multm_ps9;
  wire multm_ps10;
  wire multm_ps11;
  wire multm_ps12;
  wire multm_ps13;
  wire multm_ps14;
  wire multm_ps15;
  wire multm_ps16;
  wire multm_ps17;
  wire multm_ps18;
  wire multm_ps19;
  wire multm_ps20;
  wire multm_ps21;
  wire multm_ps22;
  wire multm_ps23;
  wire multm_ps24;
  wire multm_ps25;
  wire multm_ps26;
  wire multm_ps27;
  wire multm_ps28;
  wire multm_ps29;
  wire multm_ps30;
  wire multm_ps31;
  wire multm_ps32;
  wire multm_ps33;
  wire multm_ps34;
  wire multm_ps35;
  wire multm_ps36;
  wire multm_ps37;
  wire multm_ps38;
  wire multm_ps39;
  wire multm_ps40;
  wire multm_ps41;
  wire multm_ps42;
  wire multm_ps43;
  wire multm_ps44;
  wire multm_ps45;
  wire multm_ps46;
  wire multm_ps47;
  wire multm_ps48;
  wire multm_ps49;
  wire multm_ps50;
  wire multm_ps51;
  wire multm_ps52;
  wire multm_ps53;
  wire multm_ps54;
  wire multm_ps55;
  wire multm_ps56;
  wire multm_ps57;
  wire multm_ps58;
  wire multm_ps59;
  wire multm_ps60;
  wire multm_ps61;
  wire multm_ps62;
  wire multm_ps63;
  wire multm_ps64;
  wire multm_ps65;
  wire multm_ps66;
  wire multm_ps67;
  wire multm_ps68;
  wire multm_ps69;
  wire multm_ps70;
  wire multm_ps71;
  wire multm_ps72;
  wire multm_ps73;
  wire multm_ps74;
  wire multm_ps75;
  wire multm_ps76;
  wire multm_ps77;
  wire multm_ps78;
  wire multm_ps79;
  wire multm_ps80;
  wire multm_ps81;
  wire multm_ps82;
  wire multm_ps83;
  wire multm_ps84;
  wire multm_ps85;
  wire multm_ps86;
  wire multm_ps87;
  wire multm_ps88;
  wire multm_ps89;
  wire multm_ps90;
  wire multm_ps91;
  wire multm_ps92;
  wire multm_ps93;
  wire multm_ps94;
  wire multm_ps95;
  wire multm_ps96;
  wire multm_ps97;
  wire multm_ps98;
  wire multm_ps99;
  wire multm_ps100;
  wire multm_ps101;
  wire multm_ps102;
  wire multm_ps103;
  wire multm_ps104;
  wire multm_ps105;
  wire multm_ps106;
  wire multm_ps107;
  wire multm_ps108;
  wire multm_ps109;
  wire multm_ps110;
  wire multm_ps111;
  wire multm_ps112;
  wire multm_ps113;
  wire multm_ps114;
  wire multm_ps115;
  wire multm_ps116;
  wire multm_ps117;
  wire multm_ps118;
  wire multm_ps119;
  wire multm_ps120;
  wire multm_ps121;
  wire multm_ps122;
  wire multm_ps123;
  wire multm_ps124;
  wire multm_ps125;
  wire multm_ps126;
  wire multm_ps127;
  wire multm_ps128;
  wire multm_ps129;
  wire multm_ps130;
  wire multm_ps131;
  wire multm_ps132;
  wire multm_ps133;
  wire multm_ps134;
  wire multm_ps135;
  wire multm_ps136;
  wire multm_ps137;
  wire multm_ps138;
  wire multm_ps139;
  wire multm_ps140;
  wire multm_ps141;
  wire multm_ps142;
  wire multm_ps143;
  wire multm_ps144;
  wire multm_ps145;
  wire multm_ps146;
  wire multm_ps147;
  wire multm_ps148;
  wire multm_ps149;
  wire multm_ps150;
  wire multm_ps151;
  wire multm_ps152;
  wire multm_ps153;
  wire multm_ps154;
  wire multm_ps155;
  wire multm_ps156;
  wire multm_ps157;
  wire multm_ps158;
  wire multm_ps159;
  wire multm_ps160;
  wire multm_ps161;
  wire multm_ps162;
  wire multm_ps163;
  wire multm_ps164;
  wire multm_ps165;
  wire multm_ps166;
  wire multm_ps167;
  wire multm_ps168;
  wire multm_ps169;
  wire multm_ps170;
  wire multm_ps171;
  wire multm_ps172;
  wire multm_ps173;
  wire multm_ps174;
  wire multm_ps175;
  wire multm_ps176;
  wire multm_ps177;
  wire multm_ps178;
  wire multm_ps179;
  wire multm_ps180;
  wire multm_ps181;
  wire multm_ps182;
  wire multm_ps183;
  wire multm_ps184;
  wire multm_qcr0;
  wire multm_qcr1;
  wire multm_qcr2;
  wire multm_qcr3;
  wire multm_qcr4;
  wire multm_qcr5;
  wire multm_qcr6;
  wire multm_qcr7;
  wire multm_qcr8;
  wire multm_qcr9;
  wire multm_qcr10;
  wire multm_qcr11;
  wire multm_qcr12;
  wire multm_qcr13;
  wire multm_qcr14;
  wire multm_qcr15;
  wire multm_qcr16;
  wire multm_qcr17;
  wire multm_qcr18;
  wire multm_qcr19;
  wire multm_qcr20;
  wire multm_qcr21;
  wire multm_qcr22;
  wire multm_qcr23;
  wire multm_qcr24;
  wire multm_qcr25;
  wire multm_qcr26;
  wire multm_qcr27;
  wire multm_qcr28;
  wire multm_qcr29;
  wire multm_qcr30;
  wire multm_qcr31;
  wire multm_qcr32;
  wire multm_qcr33;
  wire multm_qcr34;
  wire multm_qcr35;
  wire multm_qcr36;
  wire multm_qcr37;
  wire multm_qcr38;
  wire multm_qcr39;
  wire multm_qcr40;
  wire multm_qcr41;
  wire multm_qcr42;
  wire multm_qcr43;
  wire multm_qcr44;
  wire multm_qcr45;
  wire multm_qcr46;
  wire multm_qcr47;
  wire multm_qcr48;
  wire multm_qcr49;
  wire multm_qcr50;
  wire multm_qcr51;
  wire multm_qcr52;
  wire multm_qcr53;
  wire multm_qcr54;
  wire multm_qcr55;
  wire multm_qcr56;
  wire multm_qcr57;
  wire multm_qcr58;
  wire multm_qcr59;
  wire multm_qcr60;
  wire multm_qcr61;
  wire multm_qcr62;
  wire multm_qcr63;
  wire multm_qcr64;
  wire multm_qcr65;
  wire multm_qcr66;
  wire multm_qcr67;
  wire multm_qcr68;
  wire multm_qcr69;
  wire multm_qcr70;
  wire multm_qcr71;
  wire multm_qcr72;
  wire multm_qcr73;
  wire multm_qcr74;
  wire multm_qcr75;
  wire multm_qcr76;
  wire multm_qcr77;
  wire multm_qcr78;
  wire multm_qcr79;
  wire multm_qcr80;
  wire multm_qcr81;
  wire multm_qcr82;
  wire multm_qcr83;
  wire multm_qcr84;
  wire multm_qcr85;
  wire multm_qcr86;
  wire multm_qcr87;
  wire multm_qcr88;
  wire multm_qcr89;
  wire multm_qcr90;
  wire multm_qcr91;
  wire multm_qcr92;
  wire multm_qcr93;
  wire multm_qcr94;
  wire multm_qcr95;
  wire multm_qcr96;
  wire multm_qcr97;
  wire multm_qcr98;
  wire multm_qcr99;
  wire multm_qcr100;
  wire multm_qcr101;
  wire multm_qcr102;
  wire multm_qcr103;
  wire multm_qcr104;
  wire multm_qcr105;
  wire multm_qcr106;
  wire multm_qcr107;
  wire multm_qcr108;
  wire multm_qcr109;
  wire multm_qcr110;
  wire multm_qcr111;
  wire multm_qcr112;
  wire multm_qcr113;
  wire multm_qcr114;
  wire multm_qcr115;
  wire multm_qcr116;
  wire multm_qcr117;
  wire multm_qcr118;
  wire multm_qcr119;
  wire multm_qcr120;
  wire multm_qcr121;
  wire multm_qcr122;
  wire multm_qcr123;
  wire multm_qcr124;
  wire multm_qcr125;
  wire multm_qcr126;
  wire multm_qcr127;
  wire multm_qcr128;
  wire multm_qcr129;
  wire multm_qcr130;
  wire multm_qcr131;
  wire multm_qcr132;
  wire multm_qcr133;
  wire multm_qcr134;
  wire multm_qcr135;
  wire multm_qcr136;
  wire multm_qcr137;
  wire multm_qcr138;
  wire multm_qcr139;
  wire multm_qcr140;
  wire multm_qcr141;
  wire multm_qcr142;
  wire multm_qcr143;
  wire multm_qcr144;
  wire multm_qcr145;
  wire multm_qcr146;
  wire multm_qcr147;
  wire multm_qcr148;
  wire multm_qcr149;
  wire multm_qcr150;
  wire multm_qcr151;
  wire multm_qcr152;
  wire multm_qcr153;
  wire multm_qcr154;
  wire multm_qcr155;
  wire multm_qcr156;
  wire multm_qcr157;
  wire multm_qcr158;
  wire multm_qcr159;
  wire multm_qcr160;
  wire multm_qcr161;
  wire multm_qcr162;
  wire multm_qcr163;
  wire multm_qcr164;
  wire multm_qcr165;
  wire multm_qcr166;
  wire multm_qcr167;
  wire multm_qcr168;
  wire multm_qcr169;
  wire multm_qcr170;
  wire multm_qcr171;
  wire multm_qcr172;
  wire multm_qcr173;
  wire multm_qcr174;
  wire multm_qcr175;
  wire multm_qcr176;
  wire multm_qcr177;
  wire multm_qcr178;
  wire multm_qcr179;
  wire multm_qcr180;
  wire multm_qcr181;
  wire multm_qcr182;
  wire multm_qcr183;
  wire multm_qcr184;
  wire multm_qsr0;
  wire multm_qsr1;
  wire multm_qsr2;
  wire multm_qsr3;
  wire multm_qsr4;
  wire multm_qsr5;
  wire multm_qsr6;
  wire multm_qsr7;
  wire multm_qsr8;
  wire multm_qsr9;
  wire multm_qsr10;
  wire multm_qsr11;
  wire multm_qsr12;
  wire multm_qsr13;
  wire multm_qsr14;
  wire multm_qsr15;
  wire multm_qsr16;
  wire multm_qsr17;
  wire multm_qsr18;
  wire multm_qsr19;
  wire multm_qsr20;
  wire multm_qsr21;
  wire multm_qsr22;
  wire multm_qsr23;
  wire multm_qsr24;
  wire multm_qsr25;
  wire multm_qsr26;
  wire multm_qsr27;
  wire multm_qsr28;
  wire multm_qsr29;
  wire multm_qsr30;
  wire multm_qsr31;
  wire multm_qsr32;
  wire multm_qsr33;
  wire multm_qsr34;
  wire multm_qsr35;
  wire multm_qsr36;
  wire multm_qsr37;
  wire multm_qsr38;
  wire multm_qsr39;
  wire multm_qsr40;
  wire multm_qsr41;
  wire multm_qsr42;
  wire multm_qsr43;
  wire multm_qsr44;
  wire multm_qsr45;
  wire multm_qsr46;
  wire multm_qsr47;
  wire multm_qsr48;
  wire multm_qsr49;
  wire multm_qsr50;
  wire multm_qsr51;
  wire multm_qsr52;
  wire multm_qsr53;
  wire multm_qsr54;
  wire multm_qsr55;
  wire multm_qsr56;
  wire multm_qsr57;
  wire multm_qsr58;
  wire multm_qsr59;
  wire multm_qsr60;
  wire multm_qsr61;
  wire multm_qsr62;
  wire multm_qsr63;
  wire multm_qsr64;
  wire multm_qsr65;
  wire multm_qsr66;
  wire multm_qsr67;
  wire multm_qsr68;
  wire multm_qsr69;
  wire multm_qsr70;
  wire multm_qsr71;
  wire multm_qsr72;
  wire multm_qsr73;
  wire multm_qsr74;
  wire multm_qsr75;
  wire multm_qsr76;
  wire multm_qsr77;
  wire multm_qsr78;
  wire multm_qsr79;
  wire multm_qsr80;
  wire multm_qsr81;
  wire multm_qsr82;
  wire multm_qsr83;
  wire multm_qsr84;
  wire multm_qsr85;
  wire multm_qsr86;
  wire multm_qsr87;
  wire multm_qsr88;
  wire multm_qsr89;
  wire multm_qsr90;
  wire multm_qsr91;
  wire multm_qsr92;
  wire multm_qsr93;
  wire multm_qsr94;
  wire multm_qsr95;
  wire multm_qsr96;
  wire multm_qsr97;
  wire multm_qsr98;
  wire multm_qsr99;
  wire multm_qsr100;
  wire multm_qsr101;
  wire multm_qsr102;
  wire multm_qsr103;
  wire multm_qsr104;
  wire multm_qsr105;
  wire multm_qsr106;
  wire multm_qsr107;
  wire multm_qsr108;
  wire multm_qsr109;
  wire multm_qsr110;
  wire multm_qsr111;
  wire multm_qsr112;
  wire multm_qsr113;
  wire multm_qsr114;
  wire multm_qsr115;
  wire multm_qsr116;
  wire multm_qsr117;
  wire multm_qsr118;
  wire multm_qsr119;
  wire multm_qsr120;
  wire multm_qsr121;
  wire multm_qsr122;
  wire multm_qsr123;
  wire multm_qsr124;
  wire multm_qsr125;
  wire multm_qsr126;
  wire multm_qsr127;
  wire multm_qsr128;
  wire multm_qsr129;
  wire multm_qsr130;
  wire multm_qsr131;
  wire multm_qsr132;
  wire multm_qsr133;
  wire multm_qsr134;
  wire multm_qsr135;
  wire multm_qsr136;
  wire multm_qsr137;
  wire multm_qsr138;
  wire multm_qsr139;
  wire multm_qsr140;
  wire multm_qsr141;
  wire multm_qsr142;
  wire multm_qsr143;
  wire multm_qsr144;
  wire multm_qsr145;
  wire multm_qsr146;
  wire multm_qsr147;
  wire multm_qsr148;
  wire multm_qsr149;
  wire multm_qsr150;
  wire multm_qsr151;
  wire multm_qsr152;
  wire multm_qsr153;
  wire multm_qsr154;
  wire multm_qsr155;
  wire multm_qsr156;
  wire multm_qsr157;
  wire multm_qsr158;
  wire multm_qsr159;
  wire multm_qsr160;
  wire multm_qsr161;
  wire multm_qsr162;
  wire multm_qsr163;
  wire multm_qsr164;
  wire multm_qsr165;
  wire multm_qsr166;
  wire multm_qsr167;
  wire multm_qsr168;
  wire multm_qsr169;
  wire multm_qsr170;
  wire multm_qsr171;
  wire multm_qsr172;
  wire multm_qsr173;
  wire multm_qsr174;
  wire multm_qsr175;
  wire multm_qsr176;
  wire multm_qsr177;
  wire multm_qsr178;
  wire multm_qsr179;
  wire multm_qsr180;
  wire multm_qsr181;
  wire multm_qsr182;
  wire multm_qsr183;
  wire multm_qsr184;
  wire multm_reduce_add3_maj3_or3_wx;
  wire multm_reduce_add3_maj3_wx;
  wire multm_reduce_add3_maj3_wy;
  wire multm_reduce_add3_maj3_xy;
  wire multm_reduce_add3_xor3_wx;
  wire multm_reduce_add3b0_maj3b_or3b_wx0;
  wire multm_reduce_add3b0_maj3b_or3b_wx1;
  wire multm_reduce_add3b0_maj3b_or3b_wx2;
  wire multm_reduce_add3b0_maj3b_or3b_wx3;
  wire multm_reduce_add3b0_maj3b_or3b_wx4;
  wire multm_reduce_add3b0_maj3b_or3b_wx5;
  wire multm_reduce_add3b0_maj3b_or3b_wx6;
  wire multm_reduce_add3b0_maj3b_or3b_wx7;
  wire multm_reduce_add3b0_maj3b_or3b_wx8;
  wire multm_reduce_add3b0_maj3b_or3b_wx9;
  wire multm_reduce_add3b0_maj3b_or3b_wx10;
  wire multm_reduce_add3b0_maj3b_or3b_wx11;
  wire multm_reduce_add3b0_maj3b_or3b_wx12;
  wire multm_reduce_add3b0_maj3b_or3b_wx13;
  wire multm_reduce_add3b0_maj3b_or3b_wx14;
  wire multm_reduce_add3b0_maj3b_or3b_wx15;
  wire multm_reduce_add3b0_maj3b_or3b_wx16;
  wire multm_reduce_add3b0_maj3b_or3b_wx17;
  wire multm_reduce_add3b0_maj3b_or3b_wx18;
  wire multm_reduce_add3b0_maj3b_or3b_wx19;
  wire multm_reduce_add3b0_maj3b_or3b_wx20;
  wire multm_reduce_add3b0_maj3b_or3b_wx21;
  wire multm_reduce_add3b0_maj3b_or3b_wx22;
  wire multm_reduce_add3b0_maj3b_or3b_wx23;
  wire multm_reduce_add3b0_maj3b_or3b_wx24;
  wire multm_reduce_add3b0_maj3b_or3b_wx25;
  wire multm_reduce_add3b0_maj3b_or3b_wx26;
  wire multm_reduce_add3b0_maj3b_or3b_wx27;
  wire multm_reduce_add3b0_maj3b_or3b_wx28;
  wire multm_reduce_add3b0_maj3b_or3b_wx29;
  wire multm_reduce_add3b0_maj3b_or3b_wx30;
  wire multm_reduce_add3b0_maj3b_or3b_wx31;
  wire multm_reduce_add3b0_maj3b_or3b_wx32;
  wire multm_reduce_add3b0_maj3b_or3b_wx33;
  wire multm_reduce_add3b0_maj3b_or3b_wx34;
  wire multm_reduce_add3b0_maj3b_or3b_wx35;
  wire multm_reduce_add3b0_maj3b_or3b_wx36;
  wire multm_reduce_add3b0_maj3b_or3b_wx37;
  wire multm_reduce_add3b0_maj3b_or3b_wx38;
  wire multm_reduce_add3b0_maj3b_or3b_wx39;
  wire multm_reduce_add3b0_maj3b_or3b_wx40;
  wire multm_reduce_add3b0_maj3b_or3b_wx41;
  wire multm_reduce_add3b0_maj3b_or3b_wx42;
  wire multm_reduce_add3b0_maj3b_or3b_wx43;
  wire multm_reduce_add3b0_maj3b_or3b_wx44;
  wire multm_reduce_add3b0_maj3b_or3b_wx45;
  wire multm_reduce_add3b0_maj3b_or3b_wx46;
  wire multm_reduce_add3b0_maj3b_or3b_wx47;
  wire multm_reduce_add3b0_maj3b_or3b_wx48;
  wire multm_reduce_add3b0_maj3b_or3b_wx49;
  wire multm_reduce_add3b0_maj3b_or3b_wx50;
  wire multm_reduce_add3b0_maj3b_or3b_wx51;
  wire multm_reduce_add3b0_maj3b_or3b_wx52;
  wire multm_reduce_add3b0_maj3b_or3b_wx53;
  wire multm_reduce_add3b0_maj3b_or3b_wx54;
  wire multm_reduce_add3b0_maj3b_or3b_wx55;
  wire multm_reduce_add3b0_maj3b_or3b_wx56;
  wire multm_reduce_add3b0_maj3b_or3b_wx57;
  wire multm_reduce_add3b0_maj3b_or3b_wx58;
  wire multm_reduce_add3b0_maj3b_or3b_wx59;
  wire multm_reduce_add3b0_maj3b_or3b_wx60;
  wire multm_reduce_add3b0_maj3b_or3b_wx61;
  wire multm_reduce_add3b0_maj3b_or3b_wx62;
  wire multm_reduce_add3b0_maj3b_or3b_wx63;
  wire multm_reduce_add3b0_maj3b_or3b_wx64;
  wire multm_reduce_add3b0_maj3b_or3b_wx65;
  wire multm_reduce_add3b0_maj3b_or3b_wx66;
  wire multm_reduce_add3b0_maj3b_or3b_wx67;
  wire multm_reduce_add3b0_maj3b_or3b_wx68;
  wire multm_reduce_add3b0_maj3b_or3b_wx69;
  wire multm_reduce_add3b0_maj3b_or3b_wx70;
  wire multm_reduce_add3b0_maj3b_or3b_wx71;
  wire multm_reduce_add3b0_maj3b_or3b_wx72;
  wire multm_reduce_add3b0_maj3b_or3b_wx73;
  wire multm_reduce_add3b0_maj3b_or3b_wx74;
  wire multm_reduce_add3b0_maj3b_or3b_wx75;
  wire multm_reduce_add3b0_maj3b_or3b_wx76;
  wire multm_reduce_add3b0_maj3b_or3b_wx77;
  wire multm_reduce_add3b0_maj3b_or3b_wx78;
  wire multm_reduce_add3b0_maj3b_or3b_wx79;
  wire multm_reduce_add3b0_maj3b_or3b_wx80;
  wire multm_reduce_add3b0_maj3b_or3b_wx81;
  wire multm_reduce_add3b0_maj3b_or3b_wx82;
  wire multm_reduce_add3b0_maj3b_or3b_wx83;
  wire multm_reduce_add3b0_maj3b_or3b_wx84;
  wire multm_reduce_add3b0_maj3b_or3b_wx85;
  wire multm_reduce_add3b0_maj3b_or3b_wx86;
  wire multm_reduce_add3b0_maj3b_or3b_wx87;
  wire multm_reduce_add3b0_maj3b_or3b_wx88;
  wire multm_reduce_add3b0_maj3b_or3b_wx89;
  wire multm_reduce_add3b0_maj3b_or3b_wx90;
  wire multm_reduce_add3b0_maj3b_or3b_wx91;
  wire multm_reduce_add3b0_maj3b_or3b_wx92;
  wire multm_reduce_add3b0_maj3b_or3b_wx93;
  wire multm_reduce_add3b0_maj3b_or3b_wx94;
  wire multm_reduce_add3b0_maj3b_or3b_wx95;
  wire multm_reduce_add3b0_maj3b_or3b_wx96;
  wire multm_reduce_add3b0_maj3b_or3b_wx97;
  wire multm_reduce_add3b0_maj3b_or3b_wx98;
  wire multm_reduce_add3b0_maj3b_or3b_wx99;
  wire multm_reduce_add3b0_maj3b_or3b_wx100;
  wire multm_reduce_add3b0_maj3b_or3b_wx101;
  wire multm_reduce_add3b0_maj3b_or3b_wx102;
  wire multm_reduce_add3b0_maj3b_or3b_wx103;
  wire multm_reduce_add3b0_maj3b_or3b_wx104;
  wire multm_reduce_add3b0_maj3b_or3b_wx105;
  wire multm_reduce_add3b0_maj3b_or3b_wx106;
  wire multm_reduce_add3b0_maj3b_or3b_wx107;
  wire multm_reduce_add3b0_maj3b_or3b_wx108;
  wire multm_reduce_add3b0_maj3b_or3b_wx109;
  wire multm_reduce_add3b0_maj3b_or3b_wx110;
  wire multm_reduce_add3b0_maj3b_or3b_wx111;
  wire multm_reduce_add3b0_maj3b_or3b_wx112;
  wire multm_reduce_add3b0_maj3b_or3b_wx113;
  wire multm_reduce_add3b0_maj3b_or3b_wx114;
  wire multm_reduce_add3b0_maj3b_or3b_wx115;
  wire multm_reduce_add3b0_maj3b_or3b_wx116;
  wire multm_reduce_add3b0_maj3b_or3b_wx117;
  wire multm_reduce_add3b0_maj3b_or3b_wx118;
  wire multm_reduce_add3b0_maj3b_or3b_wx119;
  wire multm_reduce_add3b0_maj3b_or3b_wx120;
  wire multm_reduce_add3b0_maj3b_or3b_wx121;
  wire multm_reduce_add3b0_maj3b_or3b_wx122;
  wire multm_reduce_add3b0_maj3b_or3b_wx123;
  wire multm_reduce_add3b0_maj3b_or3b_wx124;
  wire multm_reduce_add3b0_maj3b_or3b_wx125;
  wire multm_reduce_add3b0_maj3b_or3b_wx126;
  wire multm_reduce_add3b0_maj3b_or3b_wx127;
  wire multm_reduce_add3b0_maj3b_or3b_wx128;
  wire multm_reduce_add3b0_maj3b_or3b_wx129;
  wire multm_reduce_add3b0_maj3b_or3b_wx130;
  wire multm_reduce_add3b0_maj3b_or3b_wx131;
  wire multm_reduce_add3b0_maj3b_or3b_wx132;
  wire multm_reduce_add3b0_maj3b_or3b_wx133;
  wire multm_reduce_add3b0_maj3b_or3b_wx134;
  wire multm_reduce_add3b0_maj3b_or3b_wx135;
  wire multm_reduce_add3b0_maj3b_or3b_wx136;
  wire multm_reduce_add3b0_maj3b_or3b_wx137;
  wire multm_reduce_add3b0_maj3b_or3b_wx138;
  wire multm_reduce_add3b0_maj3b_or3b_wx139;
  wire multm_reduce_add3b0_maj3b_or3b_wx140;
  wire multm_reduce_add3b0_maj3b_or3b_wx141;
  wire multm_reduce_add3b0_maj3b_or3b_wx142;
  wire multm_reduce_add3b0_maj3b_or3b_wx143;
  wire multm_reduce_add3b0_maj3b_or3b_wx144;
  wire multm_reduce_add3b0_maj3b_or3b_wx145;
  wire multm_reduce_add3b0_maj3b_or3b_wx146;
  wire multm_reduce_add3b0_maj3b_or3b_wx147;
  wire multm_reduce_add3b0_maj3b_or3b_wx148;
  wire multm_reduce_add3b0_maj3b_or3b_wx149;
  wire multm_reduce_add3b0_maj3b_or3b_wx150;
  wire multm_reduce_add3b0_maj3b_or3b_wx151;
  wire multm_reduce_add3b0_maj3b_or3b_wx152;
  wire multm_reduce_add3b0_maj3b_or3b_wx153;
  wire multm_reduce_add3b0_maj3b_or3b_wx154;
  wire multm_reduce_add3b0_maj3b_or3b_wx155;
  wire multm_reduce_add3b0_maj3b_or3b_wx156;
  wire multm_reduce_add3b0_maj3b_or3b_wx157;
  wire multm_reduce_add3b0_maj3b_or3b_wx158;
  wire multm_reduce_add3b0_maj3b_or3b_wx159;
  wire multm_reduce_add3b0_maj3b_or3b_wx160;
  wire multm_reduce_add3b0_maj3b_or3b_wx161;
  wire multm_reduce_add3b0_maj3b_or3b_wx162;
  wire multm_reduce_add3b0_maj3b_or3b_wx163;
  wire multm_reduce_add3b0_maj3b_or3b_wx164;
  wire multm_reduce_add3b0_maj3b_or3b_wx165;
  wire multm_reduce_add3b0_maj3b_or3b_wx166;
  wire multm_reduce_add3b0_maj3b_or3b_wx167;
  wire multm_reduce_add3b0_maj3b_or3b_wx168;
  wire multm_reduce_add3b0_maj3b_or3b_wx169;
  wire multm_reduce_add3b0_maj3b_or3b_wx170;
  wire multm_reduce_add3b0_maj3b_or3b_wx171;
  wire multm_reduce_add3b0_maj3b_or3b_wx172;
  wire multm_reduce_add3b0_maj3b_or3b_wx173;
  wire multm_reduce_add3b0_maj3b_or3b_wx174;
  wire multm_reduce_add3b0_maj3b_or3b_wx175;
  wire multm_reduce_add3b0_maj3b_or3b_wx176;
  wire multm_reduce_add3b0_maj3b_or3b_wx177;
  wire multm_reduce_add3b0_maj3b_or3b_wx178;
  wire multm_reduce_add3b0_maj3b_or3b_wx179;
  wire multm_reduce_add3b0_maj3b_or3b_wx180;
  wire multm_reduce_add3b0_maj3b_or3b_wx181;
  wire multm_reduce_add3b0_maj3b_or3b_wx182;
  wire multm_reduce_add3b0_maj3b_wx0;
  wire multm_reduce_add3b0_maj3b_wx1;
  wire multm_reduce_add3b0_maj3b_wx2;
  wire multm_reduce_add3b0_maj3b_wx3;
  wire multm_reduce_add3b0_maj3b_wx4;
  wire multm_reduce_add3b0_maj3b_wx5;
  wire multm_reduce_add3b0_maj3b_wx6;
  wire multm_reduce_add3b0_maj3b_wx7;
  wire multm_reduce_add3b0_maj3b_wx8;
  wire multm_reduce_add3b0_maj3b_wx9;
  wire multm_reduce_add3b0_maj3b_wx10;
  wire multm_reduce_add3b0_maj3b_wx11;
  wire multm_reduce_add3b0_maj3b_wx12;
  wire multm_reduce_add3b0_maj3b_wx13;
  wire multm_reduce_add3b0_maj3b_wx14;
  wire multm_reduce_add3b0_maj3b_wx15;
  wire multm_reduce_add3b0_maj3b_wx16;
  wire multm_reduce_add3b0_maj3b_wx17;
  wire multm_reduce_add3b0_maj3b_wx18;
  wire multm_reduce_add3b0_maj3b_wx19;
  wire multm_reduce_add3b0_maj3b_wx20;
  wire multm_reduce_add3b0_maj3b_wx21;
  wire multm_reduce_add3b0_maj3b_wx22;
  wire multm_reduce_add3b0_maj3b_wx23;
  wire multm_reduce_add3b0_maj3b_wx24;
  wire multm_reduce_add3b0_maj3b_wx25;
  wire multm_reduce_add3b0_maj3b_wx26;
  wire multm_reduce_add3b0_maj3b_wx27;
  wire multm_reduce_add3b0_maj3b_wx28;
  wire multm_reduce_add3b0_maj3b_wx29;
  wire multm_reduce_add3b0_maj3b_wx30;
  wire multm_reduce_add3b0_maj3b_wx31;
  wire multm_reduce_add3b0_maj3b_wx32;
  wire multm_reduce_add3b0_maj3b_wx33;
  wire multm_reduce_add3b0_maj3b_wx34;
  wire multm_reduce_add3b0_maj3b_wx35;
  wire multm_reduce_add3b0_maj3b_wx36;
  wire multm_reduce_add3b0_maj3b_wx37;
  wire multm_reduce_add3b0_maj3b_wx38;
  wire multm_reduce_add3b0_maj3b_wx39;
  wire multm_reduce_add3b0_maj3b_wx40;
  wire multm_reduce_add3b0_maj3b_wx41;
  wire multm_reduce_add3b0_maj3b_wx42;
  wire multm_reduce_add3b0_maj3b_wx43;
  wire multm_reduce_add3b0_maj3b_wx44;
  wire multm_reduce_add3b0_maj3b_wx45;
  wire multm_reduce_add3b0_maj3b_wx46;
  wire multm_reduce_add3b0_maj3b_wx47;
  wire multm_reduce_add3b0_maj3b_wx48;
  wire multm_reduce_add3b0_maj3b_wx49;
  wire multm_reduce_add3b0_maj3b_wx50;
  wire multm_reduce_add3b0_maj3b_wx51;
  wire multm_reduce_add3b0_maj3b_wx52;
  wire multm_reduce_add3b0_maj3b_wx53;
  wire multm_reduce_add3b0_maj3b_wx54;
  wire multm_reduce_add3b0_maj3b_wx55;
  wire multm_reduce_add3b0_maj3b_wx56;
  wire multm_reduce_add3b0_maj3b_wx57;
  wire multm_reduce_add3b0_maj3b_wx58;
  wire multm_reduce_add3b0_maj3b_wx59;
  wire multm_reduce_add3b0_maj3b_wx60;
  wire multm_reduce_add3b0_maj3b_wx61;
  wire multm_reduce_add3b0_maj3b_wx62;
  wire multm_reduce_add3b0_maj3b_wx63;
  wire multm_reduce_add3b0_maj3b_wx64;
  wire multm_reduce_add3b0_maj3b_wx65;
  wire multm_reduce_add3b0_maj3b_wx66;
  wire multm_reduce_add3b0_maj3b_wx67;
  wire multm_reduce_add3b0_maj3b_wx68;
  wire multm_reduce_add3b0_maj3b_wx69;
  wire multm_reduce_add3b0_maj3b_wx70;
  wire multm_reduce_add3b0_maj3b_wx71;
  wire multm_reduce_add3b0_maj3b_wx72;
  wire multm_reduce_add3b0_maj3b_wx73;
  wire multm_reduce_add3b0_maj3b_wx74;
  wire multm_reduce_add3b0_maj3b_wx75;
  wire multm_reduce_add3b0_maj3b_wx76;
  wire multm_reduce_add3b0_maj3b_wx77;
  wire multm_reduce_add3b0_maj3b_wx78;
  wire multm_reduce_add3b0_maj3b_wx79;
  wire multm_reduce_add3b0_maj3b_wx80;
  wire multm_reduce_add3b0_maj3b_wx81;
  wire multm_reduce_add3b0_maj3b_wx82;
  wire multm_reduce_add3b0_maj3b_wx83;
  wire multm_reduce_add3b0_maj3b_wx84;
  wire multm_reduce_add3b0_maj3b_wx85;
  wire multm_reduce_add3b0_maj3b_wx86;
  wire multm_reduce_add3b0_maj3b_wx87;
  wire multm_reduce_add3b0_maj3b_wx88;
  wire multm_reduce_add3b0_maj3b_wx89;
  wire multm_reduce_add3b0_maj3b_wx90;
  wire multm_reduce_add3b0_maj3b_wx91;
  wire multm_reduce_add3b0_maj3b_wx92;
  wire multm_reduce_add3b0_maj3b_wx93;
  wire multm_reduce_add3b0_maj3b_wx94;
  wire multm_reduce_add3b0_maj3b_wx95;
  wire multm_reduce_add3b0_maj3b_wx96;
  wire multm_reduce_add3b0_maj3b_wx97;
  wire multm_reduce_add3b0_maj3b_wx98;
  wire multm_reduce_add3b0_maj3b_wx99;
  wire multm_reduce_add3b0_maj3b_wx100;
  wire multm_reduce_add3b0_maj3b_wx101;
  wire multm_reduce_add3b0_maj3b_wx102;
  wire multm_reduce_add3b0_maj3b_wx103;
  wire multm_reduce_add3b0_maj3b_wx104;
  wire multm_reduce_add3b0_maj3b_wx105;
  wire multm_reduce_add3b0_maj3b_wx106;
  wire multm_reduce_add3b0_maj3b_wx107;
  wire multm_reduce_add3b0_maj3b_wx108;
  wire multm_reduce_add3b0_maj3b_wx109;
  wire multm_reduce_add3b0_maj3b_wx110;
  wire multm_reduce_add3b0_maj3b_wx111;
  wire multm_reduce_add3b0_maj3b_wx112;
  wire multm_reduce_add3b0_maj3b_wx113;
  wire multm_reduce_add3b0_maj3b_wx114;
  wire multm_reduce_add3b0_maj3b_wx115;
  wire multm_reduce_add3b0_maj3b_wx116;
  wire multm_reduce_add3b0_maj3b_wx117;
  wire multm_reduce_add3b0_maj3b_wx118;
  wire multm_reduce_add3b0_maj3b_wx119;
  wire multm_reduce_add3b0_maj3b_wx120;
  wire multm_reduce_add3b0_maj3b_wx121;
  wire multm_reduce_add3b0_maj3b_wx122;
  wire multm_reduce_add3b0_maj3b_wx123;
  wire multm_reduce_add3b0_maj3b_wx124;
  wire multm_reduce_add3b0_maj3b_wx125;
  wire multm_reduce_add3b0_maj3b_wx126;
  wire multm_reduce_add3b0_maj3b_wx127;
  wire multm_reduce_add3b0_maj3b_wx128;
  wire multm_reduce_add3b0_maj3b_wx129;
  wire multm_reduce_add3b0_maj3b_wx130;
  wire multm_reduce_add3b0_maj3b_wx131;
  wire multm_reduce_add3b0_maj3b_wx132;
  wire multm_reduce_add3b0_maj3b_wx133;
  wire multm_reduce_add3b0_maj3b_wx134;
  wire multm_reduce_add3b0_maj3b_wx135;
  wire multm_reduce_add3b0_maj3b_wx136;
  wire multm_reduce_add3b0_maj3b_wx137;
  wire multm_reduce_add3b0_maj3b_wx138;
  wire multm_reduce_add3b0_maj3b_wx139;
  wire multm_reduce_add3b0_maj3b_wx140;
  wire multm_reduce_add3b0_maj3b_wx141;
  wire multm_reduce_add3b0_maj3b_wx142;
  wire multm_reduce_add3b0_maj3b_wx143;
  wire multm_reduce_add3b0_maj3b_wx144;
  wire multm_reduce_add3b0_maj3b_wx145;
  wire multm_reduce_add3b0_maj3b_wx146;
  wire multm_reduce_add3b0_maj3b_wx147;
  wire multm_reduce_add3b0_maj3b_wx148;
  wire multm_reduce_add3b0_maj3b_wx149;
  wire multm_reduce_add3b0_maj3b_wx150;
  wire multm_reduce_add3b0_maj3b_wx151;
  wire multm_reduce_add3b0_maj3b_wx152;
  wire multm_reduce_add3b0_maj3b_wx153;
  wire multm_reduce_add3b0_maj3b_wx154;
  wire multm_reduce_add3b0_maj3b_wx155;
  wire multm_reduce_add3b0_maj3b_wx156;
  wire multm_reduce_add3b0_maj3b_wx157;
  wire multm_reduce_add3b0_maj3b_wx158;
  wire multm_reduce_add3b0_maj3b_wx159;
  wire multm_reduce_add3b0_maj3b_wx160;
  wire multm_reduce_add3b0_maj3b_wx161;
  wire multm_reduce_add3b0_maj3b_wx162;
  wire multm_reduce_add3b0_maj3b_wx163;
  wire multm_reduce_add3b0_maj3b_wx164;
  wire multm_reduce_add3b0_maj3b_wx165;
  wire multm_reduce_add3b0_maj3b_wx166;
  wire multm_reduce_add3b0_maj3b_wx167;
  wire multm_reduce_add3b0_maj3b_wx168;
  wire multm_reduce_add3b0_maj3b_wx169;
  wire multm_reduce_add3b0_maj3b_wx170;
  wire multm_reduce_add3b0_maj3b_wx171;
  wire multm_reduce_add3b0_maj3b_wx172;
  wire multm_reduce_add3b0_maj3b_wx173;
  wire multm_reduce_add3b0_maj3b_wx174;
  wire multm_reduce_add3b0_maj3b_wx175;
  wire multm_reduce_add3b0_maj3b_wx176;
  wire multm_reduce_add3b0_maj3b_wx177;
  wire multm_reduce_add3b0_maj3b_wx178;
  wire multm_reduce_add3b0_maj3b_wx179;
  wire multm_reduce_add3b0_maj3b_wx180;
  wire multm_reduce_add3b0_maj3b_wx181;
  wire multm_reduce_add3b0_maj3b_wx182;
  wire multm_reduce_add3b0_maj3b_wy0;
  wire multm_reduce_add3b0_maj3b_wy1;
  wire multm_reduce_add3b0_maj3b_wy2;
  wire multm_reduce_add3b0_maj3b_wy3;
  wire multm_reduce_add3b0_maj3b_wy4;
  wire multm_reduce_add3b0_maj3b_wy5;
  wire multm_reduce_add3b0_maj3b_wy6;
  wire multm_reduce_add3b0_maj3b_wy7;
  wire multm_reduce_add3b0_maj3b_wy8;
  wire multm_reduce_add3b0_maj3b_wy9;
  wire multm_reduce_add3b0_maj3b_wy10;
  wire multm_reduce_add3b0_maj3b_wy11;
  wire multm_reduce_add3b0_maj3b_wy12;
  wire multm_reduce_add3b0_maj3b_wy13;
  wire multm_reduce_add3b0_maj3b_wy14;
  wire multm_reduce_add3b0_maj3b_wy15;
  wire multm_reduce_add3b0_maj3b_wy16;
  wire multm_reduce_add3b0_maj3b_wy17;
  wire multm_reduce_add3b0_maj3b_wy18;
  wire multm_reduce_add3b0_maj3b_wy19;
  wire multm_reduce_add3b0_maj3b_wy20;
  wire multm_reduce_add3b0_maj3b_wy21;
  wire multm_reduce_add3b0_maj3b_wy22;
  wire multm_reduce_add3b0_maj3b_wy23;
  wire multm_reduce_add3b0_maj3b_wy24;
  wire multm_reduce_add3b0_maj3b_wy25;
  wire multm_reduce_add3b0_maj3b_wy26;
  wire multm_reduce_add3b0_maj3b_wy27;
  wire multm_reduce_add3b0_maj3b_wy28;
  wire multm_reduce_add3b0_maj3b_wy29;
  wire multm_reduce_add3b0_maj3b_wy30;
  wire multm_reduce_add3b0_maj3b_wy31;
  wire multm_reduce_add3b0_maj3b_wy32;
  wire multm_reduce_add3b0_maj3b_wy33;
  wire multm_reduce_add3b0_maj3b_wy34;
  wire multm_reduce_add3b0_maj3b_wy35;
  wire multm_reduce_add3b0_maj3b_wy36;
  wire multm_reduce_add3b0_maj3b_wy37;
  wire multm_reduce_add3b0_maj3b_wy38;
  wire multm_reduce_add3b0_maj3b_wy39;
  wire multm_reduce_add3b0_maj3b_wy40;
  wire multm_reduce_add3b0_maj3b_wy41;
  wire multm_reduce_add3b0_maj3b_wy42;
  wire multm_reduce_add3b0_maj3b_wy43;
  wire multm_reduce_add3b0_maj3b_wy44;
  wire multm_reduce_add3b0_maj3b_wy45;
  wire multm_reduce_add3b0_maj3b_wy46;
  wire multm_reduce_add3b0_maj3b_wy47;
  wire multm_reduce_add3b0_maj3b_wy48;
  wire multm_reduce_add3b0_maj3b_wy49;
  wire multm_reduce_add3b0_maj3b_wy50;
  wire multm_reduce_add3b0_maj3b_wy51;
  wire multm_reduce_add3b0_maj3b_wy52;
  wire multm_reduce_add3b0_maj3b_wy53;
  wire multm_reduce_add3b0_maj3b_wy54;
  wire multm_reduce_add3b0_maj3b_wy55;
  wire multm_reduce_add3b0_maj3b_wy56;
  wire multm_reduce_add3b0_maj3b_wy57;
  wire multm_reduce_add3b0_maj3b_wy58;
  wire multm_reduce_add3b0_maj3b_wy59;
  wire multm_reduce_add3b0_maj3b_wy60;
  wire multm_reduce_add3b0_maj3b_wy61;
  wire multm_reduce_add3b0_maj3b_wy62;
  wire multm_reduce_add3b0_maj3b_wy63;
  wire multm_reduce_add3b0_maj3b_wy64;
  wire multm_reduce_add3b0_maj3b_wy65;
  wire multm_reduce_add3b0_maj3b_wy66;
  wire multm_reduce_add3b0_maj3b_wy67;
  wire multm_reduce_add3b0_maj3b_wy68;
  wire multm_reduce_add3b0_maj3b_wy69;
  wire multm_reduce_add3b0_maj3b_wy70;
  wire multm_reduce_add3b0_maj3b_wy71;
  wire multm_reduce_add3b0_maj3b_wy72;
  wire multm_reduce_add3b0_maj3b_wy73;
  wire multm_reduce_add3b0_maj3b_wy74;
  wire multm_reduce_add3b0_maj3b_wy75;
  wire multm_reduce_add3b0_maj3b_wy76;
  wire multm_reduce_add3b0_maj3b_wy77;
  wire multm_reduce_add3b0_maj3b_wy78;
  wire multm_reduce_add3b0_maj3b_wy79;
  wire multm_reduce_add3b0_maj3b_wy80;
  wire multm_reduce_add3b0_maj3b_wy81;
  wire multm_reduce_add3b0_maj3b_wy82;
  wire multm_reduce_add3b0_maj3b_wy83;
  wire multm_reduce_add3b0_maj3b_wy84;
  wire multm_reduce_add3b0_maj3b_wy85;
  wire multm_reduce_add3b0_maj3b_wy86;
  wire multm_reduce_add3b0_maj3b_wy87;
  wire multm_reduce_add3b0_maj3b_wy88;
  wire multm_reduce_add3b0_maj3b_wy89;
  wire multm_reduce_add3b0_maj3b_wy90;
  wire multm_reduce_add3b0_maj3b_wy91;
  wire multm_reduce_add3b0_maj3b_wy92;
  wire multm_reduce_add3b0_maj3b_wy93;
  wire multm_reduce_add3b0_maj3b_wy94;
  wire multm_reduce_add3b0_maj3b_wy95;
  wire multm_reduce_add3b0_maj3b_wy96;
  wire multm_reduce_add3b0_maj3b_wy97;
  wire multm_reduce_add3b0_maj3b_wy98;
  wire multm_reduce_add3b0_maj3b_wy99;
  wire multm_reduce_add3b0_maj3b_wy100;
  wire multm_reduce_add3b0_maj3b_wy101;
  wire multm_reduce_add3b0_maj3b_wy102;
  wire multm_reduce_add3b0_maj3b_wy103;
  wire multm_reduce_add3b0_maj3b_wy104;
  wire multm_reduce_add3b0_maj3b_wy105;
  wire multm_reduce_add3b0_maj3b_wy106;
  wire multm_reduce_add3b0_maj3b_wy107;
  wire multm_reduce_add3b0_maj3b_wy108;
  wire multm_reduce_add3b0_maj3b_wy109;
  wire multm_reduce_add3b0_maj3b_wy110;
  wire multm_reduce_add3b0_maj3b_wy111;
  wire multm_reduce_add3b0_maj3b_wy112;
  wire multm_reduce_add3b0_maj3b_wy113;
  wire multm_reduce_add3b0_maj3b_wy114;
  wire multm_reduce_add3b0_maj3b_wy115;
  wire multm_reduce_add3b0_maj3b_wy116;
  wire multm_reduce_add3b0_maj3b_wy117;
  wire multm_reduce_add3b0_maj3b_wy118;
  wire multm_reduce_add3b0_maj3b_wy119;
  wire multm_reduce_add3b0_maj3b_wy120;
  wire multm_reduce_add3b0_maj3b_wy121;
  wire multm_reduce_add3b0_maj3b_wy122;
  wire multm_reduce_add3b0_maj3b_wy123;
  wire multm_reduce_add3b0_maj3b_wy124;
  wire multm_reduce_add3b0_maj3b_wy125;
  wire multm_reduce_add3b0_maj3b_wy126;
  wire multm_reduce_add3b0_maj3b_wy127;
  wire multm_reduce_add3b0_maj3b_wy128;
  wire multm_reduce_add3b0_maj3b_wy129;
  wire multm_reduce_add3b0_maj3b_wy130;
  wire multm_reduce_add3b0_maj3b_wy131;
  wire multm_reduce_add3b0_maj3b_wy132;
  wire multm_reduce_add3b0_maj3b_wy133;
  wire multm_reduce_add3b0_maj3b_wy134;
  wire multm_reduce_add3b0_maj3b_wy135;
  wire multm_reduce_add3b0_maj3b_wy136;
  wire multm_reduce_add3b0_maj3b_wy137;
  wire multm_reduce_add3b0_maj3b_wy138;
  wire multm_reduce_add3b0_maj3b_wy139;
  wire multm_reduce_add3b0_maj3b_wy140;
  wire multm_reduce_add3b0_maj3b_wy141;
  wire multm_reduce_add3b0_maj3b_wy142;
  wire multm_reduce_add3b0_maj3b_wy143;
  wire multm_reduce_add3b0_maj3b_wy144;
  wire multm_reduce_add3b0_maj3b_wy145;
  wire multm_reduce_add3b0_maj3b_wy146;
  wire multm_reduce_add3b0_maj3b_wy147;
  wire multm_reduce_add3b0_maj3b_wy148;
  wire multm_reduce_add3b0_maj3b_wy149;
  wire multm_reduce_add3b0_maj3b_wy150;
  wire multm_reduce_add3b0_maj3b_wy151;
  wire multm_reduce_add3b0_maj3b_wy152;
  wire multm_reduce_add3b0_maj3b_wy153;
  wire multm_reduce_add3b0_maj3b_wy154;
  wire multm_reduce_add3b0_maj3b_wy155;
  wire multm_reduce_add3b0_maj3b_wy156;
  wire multm_reduce_add3b0_maj3b_wy157;
  wire multm_reduce_add3b0_maj3b_wy158;
  wire multm_reduce_add3b0_maj3b_wy159;
  wire multm_reduce_add3b0_maj3b_wy160;
  wire multm_reduce_add3b0_maj3b_wy161;
  wire multm_reduce_add3b0_maj3b_wy162;
  wire multm_reduce_add3b0_maj3b_wy163;
  wire multm_reduce_add3b0_maj3b_wy164;
  wire multm_reduce_add3b0_maj3b_wy165;
  wire multm_reduce_add3b0_maj3b_wy166;
  wire multm_reduce_add3b0_maj3b_wy167;
  wire multm_reduce_add3b0_maj3b_wy168;
  wire multm_reduce_add3b0_maj3b_wy169;
  wire multm_reduce_add3b0_maj3b_wy170;
  wire multm_reduce_add3b0_maj3b_wy171;
  wire multm_reduce_add3b0_maj3b_wy172;
  wire multm_reduce_add3b0_maj3b_wy173;
  wire multm_reduce_add3b0_maj3b_wy174;
  wire multm_reduce_add3b0_maj3b_wy175;
  wire multm_reduce_add3b0_maj3b_wy176;
  wire multm_reduce_add3b0_maj3b_wy177;
  wire multm_reduce_add3b0_maj3b_wy178;
  wire multm_reduce_add3b0_maj3b_wy179;
  wire multm_reduce_add3b0_maj3b_wy180;
  wire multm_reduce_add3b0_maj3b_wy181;
  wire multm_reduce_add3b0_maj3b_wy182;
  wire multm_reduce_add3b0_maj3b_xy0;
  wire multm_reduce_add3b0_maj3b_xy1;
  wire multm_reduce_add3b0_maj3b_xy2;
  wire multm_reduce_add3b0_maj3b_xy3;
  wire multm_reduce_add3b0_maj3b_xy4;
  wire multm_reduce_add3b0_maj3b_xy5;
  wire multm_reduce_add3b0_maj3b_xy6;
  wire multm_reduce_add3b0_maj3b_xy7;
  wire multm_reduce_add3b0_maj3b_xy8;
  wire multm_reduce_add3b0_maj3b_xy9;
  wire multm_reduce_add3b0_maj3b_xy10;
  wire multm_reduce_add3b0_maj3b_xy11;
  wire multm_reduce_add3b0_maj3b_xy12;
  wire multm_reduce_add3b0_maj3b_xy13;
  wire multm_reduce_add3b0_maj3b_xy14;
  wire multm_reduce_add3b0_maj3b_xy15;
  wire multm_reduce_add3b0_maj3b_xy16;
  wire multm_reduce_add3b0_maj3b_xy17;
  wire multm_reduce_add3b0_maj3b_xy18;
  wire multm_reduce_add3b0_maj3b_xy19;
  wire multm_reduce_add3b0_maj3b_xy20;
  wire multm_reduce_add3b0_maj3b_xy21;
  wire multm_reduce_add3b0_maj3b_xy22;
  wire multm_reduce_add3b0_maj3b_xy23;
  wire multm_reduce_add3b0_maj3b_xy24;
  wire multm_reduce_add3b0_maj3b_xy25;
  wire multm_reduce_add3b0_maj3b_xy26;
  wire multm_reduce_add3b0_maj3b_xy27;
  wire multm_reduce_add3b0_maj3b_xy28;
  wire multm_reduce_add3b0_maj3b_xy29;
  wire multm_reduce_add3b0_maj3b_xy30;
  wire multm_reduce_add3b0_maj3b_xy31;
  wire multm_reduce_add3b0_maj3b_xy32;
  wire multm_reduce_add3b0_maj3b_xy33;
  wire multm_reduce_add3b0_maj3b_xy34;
  wire multm_reduce_add3b0_maj3b_xy35;
  wire multm_reduce_add3b0_maj3b_xy36;
  wire multm_reduce_add3b0_maj3b_xy37;
  wire multm_reduce_add3b0_maj3b_xy38;
  wire multm_reduce_add3b0_maj3b_xy39;
  wire multm_reduce_add3b0_maj3b_xy40;
  wire multm_reduce_add3b0_maj3b_xy41;
  wire multm_reduce_add3b0_maj3b_xy42;
  wire multm_reduce_add3b0_maj3b_xy43;
  wire multm_reduce_add3b0_maj3b_xy44;
  wire multm_reduce_add3b0_maj3b_xy45;
  wire multm_reduce_add3b0_maj3b_xy46;
  wire multm_reduce_add3b0_maj3b_xy47;
  wire multm_reduce_add3b0_maj3b_xy48;
  wire multm_reduce_add3b0_maj3b_xy49;
  wire multm_reduce_add3b0_maj3b_xy50;
  wire multm_reduce_add3b0_maj3b_xy51;
  wire multm_reduce_add3b0_maj3b_xy52;
  wire multm_reduce_add3b0_maj3b_xy53;
  wire multm_reduce_add3b0_maj3b_xy54;
  wire multm_reduce_add3b0_maj3b_xy55;
  wire multm_reduce_add3b0_maj3b_xy56;
  wire multm_reduce_add3b0_maj3b_xy57;
  wire multm_reduce_add3b0_maj3b_xy58;
  wire multm_reduce_add3b0_maj3b_xy59;
  wire multm_reduce_add3b0_maj3b_xy60;
  wire multm_reduce_add3b0_maj3b_xy61;
  wire multm_reduce_add3b0_maj3b_xy62;
  wire multm_reduce_add3b0_maj3b_xy63;
  wire multm_reduce_add3b0_maj3b_xy64;
  wire multm_reduce_add3b0_maj3b_xy65;
  wire multm_reduce_add3b0_maj3b_xy66;
  wire multm_reduce_add3b0_maj3b_xy67;
  wire multm_reduce_add3b0_maj3b_xy68;
  wire multm_reduce_add3b0_maj3b_xy69;
  wire multm_reduce_add3b0_maj3b_xy70;
  wire multm_reduce_add3b0_maj3b_xy71;
  wire multm_reduce_add3b0_maj3b_xy72;
  wire multm_reduce_add3b0_maj3b_xy73;
  wire multm_reduce_add3b0_maj3b_xy74;
  wire multm_reduce_add3b0_maj3b_xy75;
  wire multm_reduce_add3b0_maj3b_xy76;
  wire multm_reduce_add3b0_maj3b_xy77;
  wire multm_reduce_add3b0_maj3b_xy78;
  wire multm_reduce_add3b0_maj3b_xy79;
  wire multm_reduce_add3b0_maj3b_xy80;
  wire multm_reduce_add3b0_maj3b_xy81;
  wire multm_reduce_add3b0_maj3b_xy82;
  wire multm_reduce_add3b0_maj3b_xy83;
  wire multm_reduce_add3b0_maj3b_xy84;
  wire multm_reduce_add3b0_maj3b_xy85;
  wire multm_reduce_add3b0_maj3b_xy86;
  wire multm_reduce_add3b0_maj3b_xy87;
  wire multm_reduce_add3b0_maj3b_xy88;
  wire multm_reduce_add3b0_maj3b_xy89;
  wire multm_reduce_add3b0_maj3b_xy90;
  wire multm_reduce_add3b0_maj3b_xy91;
  wire multm_reduce_add3b0_maj3b_xy92;
  wire multm_reduce_add3b0_maj3b_xy93;
  wire multm_reduce_add3b0_maj3b_xy94;
  wire multm_reduce_add3b0_maj3b_xy95;
  wire multm_reduce_add3b0_maj3b_xy96;
  wire multm_reduce_add3b0_maj3b_xy97;
  wire multm_reduce_add3b0_maj3b_xy98;
  wire multm_reduce_add3b0_maj3b_xy99;
  wire multm_reduce_add3b0_maj3b_xy100;
  wire multm_reduce_add3b0_maj3b_xy101;
  wire multm_reduce_add3b0_maj3b_xy102;
  wire multm_reduce_add3b0_maj3b_xy103;
  wire multm_reduce_add3b0_maj3b_xy104;
  wire multm_reduce_add3b0_maj3b_xy105;
  wire multm_reduce_add3b0_maj3b_xy106;
  wire multm_reduce_add3b0_maj3b_xy107;
  wire multm_reduce_add3b0_maj3b_xy108;
  wire multm_reduce_add3b0_maj3b_xy109;
  wire multm_reduce_add3b0_maj3b_xy110;
  wire multm_reduce_add3b0_maj3b_xy111;
  wire multm_reduce_add3b0_maj3b_xy112;
  wire multm_reduce_add3b0_maj3b_xy113;
  wire multm_reduce_add3b0_maj3b_xy114;
  wire multm_reduce_add3b0_maj3b_xy115;
  wire multm_reduce_add3b0_maj3b_xy116;
  wire multm_reduce_add3b0_maj3b_xy117;
  wire multm_reduce_add3b0_maj3b_xy118;
  wire multm_reduce_add3b0_maj3b_xy119;
  wire multm_reduce_add3b0_maj3b_xy120;
  wire multm_reduce_add3b0_maj3b_xy121;
  wire multm_reduce_add3b0_maj3b_xy122;
  wire multm_reduce_add3b0_maj3b_xy123;
  wire multm_reduce_add3b0_maj3b_xy124;
  wire multm_reduce_add3b0_maj3b_xy125;
  wire multm_reduce_add3b0_maj3b_xy126;
  wire multm_reduce_add3b0_maj3b_xy127;
  wire multm_reduce_add3b0_maj3b_xy128;
  wire multm_reduce_add3b0_maj3b_xy129;
  wire multm_reduce_add3b0_maj3b_xy130;
  wire multm_reduce_add3b0_maj3b_xy131;
  wire multm_reduce_add3b0_maj3b_xy132;
  wire multm_reduce_add3b0_maj3b_xy133;
  wire multm_reduce_add3b0_maj3b_xy134;
  wire multm_reduce_add3b0_maj3b_xy135;
  wire multm_reduce_add3b0_maj3b_xy136;
  wire multm_reduce_add3b0_maj3b_xy137;
  wire multm_reduce_add3b0_maj3b_xy138;
  wire multm_reduce_add3b0_maj3b_xy139;
  wire multm_reduce_add3b0_maj3b_xy140;
  wire multm_reduce_add3b0_maj3b_xy141;
  wire multm_reduce_add3b0_maj3b_xy142;
  wire multm_reduce_add3b0_maj3b_xy143;
  wire multm_reduce_add3b0_maj3b_xy144;
  wire multm_reduce_add3b0_maj3b_xy145;
  wire multm_reduce_add3b0_maj3b_xy146;
  wire multm_reduce_add3b0_maj3b_xy147;
  wire multm_reduce_add3b0_maj3b_xy148;
  wire multm_reduce_add3b0_maj3b_xy149;
  wire multm_reduce_add3b0_maj3b_xy150;
  wire multm_reduce_add3b0_maj3b_xy151;
  wire multm_reduce_add3b0_maj3b_xy152;
  wire multm_reduce_add3b0_maj3b_xy153;
  wire multm_reduce_add3b0_maj3b_xy154;
  wire multm_reduce_add3b0_maj3b_xy155;
  wire multm_reduce_add3b0_maj3b_xy156;
  wire multm_reduce_add3b0_maj3b_xy157;
  wire multm_reduce_add3b0_maj3b_xy158;
  wire multm_reduce_add3b0_maj3b_xy159;
  wire multm_reduce_add3b0_maj3b_xy160;
  wire multm_reduce_add3b0_maj3b_xy161;
  wire multm_reduce_add3b0_maj3b_xy162;
  wire multm_reduce_add3b0_maj3b_xy163;
  wire multm_reduce_add3b0_maj3b_xy164;
  wire multm_reduce_add3b0_maj3b_xy165;
  wire multm_reduce_add3b0_maj3b_xy166;
  wire multm_reduce_add3b0_maj3b_xy167;
  wire multm_reduce_add3b0_maj3b_xy168;
  wire multm_reduce_add3b0_maj3b_xy169;
  wire multm_reduce_add3b0_maj3b_xy170;
  wire multm_reduce_add3b0_maj3b_xy171;
  wire multm_reduce_add3b0_maj3b_xy172;
  wire multm_reduce_add3b0_maj3b_xy173;
  wire multm_reduce_add3b0_maj3b_xy174;
  wire multm_reduce_add3b0_maj3b_xy175;
  wire multm_reduce_add3b0_maj3b_xy176;
  wire multm_reduce_add3b0_maj3b_xy177;
  wire multm_reduce_add3b0_maj3b_xy178;
  wire multm_reduce_add3b0_maj3b_xy179;
  wire multm_reduce_add3b0_maj3b_xy180;
  wire multm_reduce_add3b0_maj3b_xy181;
  wire multm_reduce_add3b0_maj3b_xy182;
  wire multm_reduce_add3b0_xor3b_wx0;
  wire multm_reduce_add3b0_xor3b_wx1;
  wire multm_reduce_add3b0_xor3b_wx2;
  wire multm_reduce_add3b0_xor3b_wx3;
  wire multm_reduce_add3b0_xor3b_wx4;
  wire multm_reduce_add3b0_xor3b_wx5;
  wire multm_reduce_add3b0_xor3b_wx6;
  wire multm_reduce_add3b0_xor3b_wx7;
  wire multm_reduce_add3b0_xor3b_wx8;
  wire multm_reduce_add3b0_xor3b_wx9;
  wire multm_reduce_add3b0_xor3b_wx10;
  wire multm_reduce_add3b0_xor3b_wx11;
  wire multm_reduce_add3b0_xor3b_wx12;
  wire multm_reduce_add3b0_xor3b_wx13;
  wire multm_reduce_add3b0_xor3b_wx14;
  wire multm_reduce_add3b0_xor3b_wx15;
  wire multm_reduce_add3b0_xor3b_wx16;
  wire multm_reduce_add3b0_xor3b_wx17;
  wire multm_reduce_add3b0_xor3b_wx18;
  wire multm_reduce_add3b0_xor3b_wx19;
  wire multm_reduce_add3b0_xor3b_wx20;
  wire multm_reduce_add3b0_xor3b_wx21;
  wire multm_reduce_add3b0_xor3b_wx22;
  wire multm_reduce_add3b0_xor3b_wx23;
  wire multm_reduce_add3b0_xor3b_wx24;
  wire multm_reduce_add3b0_xor3b_wx25;
  wire multm_reduce_add3b0_xor3b_wx26;
  wire multm_reduce_add3b0_xor3b_wx27;
  wire multm_reduce_add3b0_xor3b_wx28;
  wire multm_reduce_add3b0_xor3b_wx29;
  wire multm_reduce_add3b0_xor3b_wx30;
  wire multm_reduce_add3b0_xor3b_wx31;
  wire multm_reduce_add3b0_xor3b_wx32;
  wire multm_reduce_add3b0_xor3b_wx33;
  wire multm_reduce_add3b0_xor3b_wx34;
  wire multm_reduce_add3b0_xor3b_wx35;
  wire multm_reduce_add3b0_xor3b_wx36;
  wire multm_reduce_add3b0_xor3b_wx37;
  wire multm_reduce_add3b0_xor3b_wx38;
  wire multm_reduce_add3b0_xor3b_wx39;
  wire multm_reduce_add3b0_xor3b_wx40;
  wire multm_reduce_add3b0_xor3b_wx41;
  wire multm_reduce_add3b0_xor3b_wx42;
  wire multm_reduce_add3b0_xor3b_wx43;
  wire multm_reduce_add3b0_xor3b_wx44;
  wire multm_reduce_add3b0_xor3b_wx45;
  wire multm_reduce_add3b0_xor3b_wx46;
  wire multm_reduce_add3b0_xor3b_wx47;
  wire multm_reduce_add3b0_xor3b_wx48;
  wire multm_reduce_add3b0_xor3b_wx49;
  wire multm_reduce_add3b0_xor3b_wx50;
  wire multm_reduce_add3b0_xor3b_wx51;
  wire multm_reduce_add3b0_xor3b_wx52;
  wire multm_reduce_add3b0_xor3b_wx53;
  wire multm_reduce_add3b0_xor3b_wx54;
  wire multm_reduce_add3b0_xor3b_wx55;
  wire multm_reduce_add3b0_xor3b_wx56;
  wire multm_reduce_add3b0_xor3b_wx57;
  wire multm_reduce_add3b0_xor3b_wx58;
  wire multm_reduce_add3b0_xor3b_wx59;
  wire multm_reduce_add3b0_xor3b_wx60;
  wire multm_reduce_add3b0_xor3b_wx61;
  wire multm_reduce_add3b0_xor3b_wx62;
  wire multm_reduce_add3b0_xor3b_wx63;
  wire multm_reduce_add3b0_xor3b_wx64;
  wire multm_reduce_add3b0_xor3b_wx65;
  wire multm_reduce_add3b0_xor3b_wx66;
  wire multm_reduce_add3b0_xor3b_wx67;
  wire multm_reduce_add3b0_xor3b_wx68;
  wire multm_reduce_add3b0_xor3b_wx69;
  wire multm_reduce_add3b0_xor3b_wx70;
  wire multm_reduce_add3b0_xor3b_wx71;
  wire multm_reduce_add3b0_xor3b_wx72;
  wire multm_reduce_add3b0_xor3b_wx73;
  wire multm_reduce_add3b0_xor3b_wx74;
  wire multm_reduce_add3b0_xor3b_wx75;
  wire multm_reduce_add3b0_xor3b_wx76;
  wire multm_reduce_add3b0_xor3b_wx77;
  wire multm_reduce_add3b0_xor3b_wx78;
  wire multm_reduce_add3b0_xor3b_wx79;
  wire multm_reduce_add3b0_xor3b_wx80;
  wire multm_reduce_add3b0_xor3b_wx81;
  wire multm_reduce_add3b0_xor3b_wx82;
  wire multm_reduce_add3b0_xor3b_wx83;
  wire multm_reduce_add3b0_xor3b_wx84;
  wire multm_reduce_add3b0_xor3b_wx85;
  wire multm_reduce_add3b0_xor3b_wx86;
  wire multm_reduce_add3b0_xor3b_wx87;
  wire multm_reduce_add3b0_xor3b_wx88;
  wire multm_reduce_add3b0_xor3b_wx89;
  wire multm_reduce_add3b0_xor3b_wx90;
  wire multm_reduce_add3b0_xor3b_wx91;
  wire multm_reduce_add3b0_xor3b_wx92;
  wire multm_reduce_add3b0_xor3b_wx93;
  wire multm_reduce_add3b0_xor3b_wx94;
  wire multm_reduce_add3b0_xor3b_wx95;
  wire multm_reduce_add3b0_xor3b_wx96;
  wire multm_reduce_add3b0_xor3b_wx97;
  wire multm_reduce_add3b0_xor3b_wx98;
  wire multm_reduce_add3b0_xor3b_wx99;
  wire multm_reduce_add3b0_xor3b_wx100;
  wire multm_reduce_add3b0_xor3b_wx101;
  wire multm_reduce_add3b0_xor3b_wx102;
  wire multm_reduce_add3b0_xor3b_wx103;
  wire multm_reduce_add3b0_xor3b_wx104;
  wire multm_reduce_add3b0_xor3b_wx105;
  wire multm_reduce_add3b0_xor3b_wx106;
  wire multm_reduce_add3b0_xor3b_wx107;
  wire multm_reduce_add3b0_xor3b_wx108;
  wire multm_reduce_add3b0_xor3b_wx109;
  wire multm_reduce_add3b0_xor3b_wx110;
  wire multm_reduce_add3b0_xor3b_wx111;
  wire multm_reduce_add3b0_xor3b_wx112;
  wire multm_reduce_add3b0_xor3b_wx113;
  wire multm_reduce_add3b0_xor3b_wx114;
  wire multm_reduce_add3b0_xor3b_wx115;
  wire multm_reduce_add3b0_xor3b_wx116;
  wire multm_reduce_add3b0_xor3b_wx117;
  wire multm_reduce_add3b0_xor3b_wx118;
  wire multm_reduce_add3b0_xor3b_wx119;
  wire multm_reduce_add3b0_xor3b_wx120;
  wire multm_reduce_add3b0_xor3b_wx121;
  wire multm_reduce_add3b0_xor3b_wx122;
  wire multm_reduce_add3b0_xor3b_wx123;
  wire multm_reduce_add3b0_xor3b_wx124;
  wire multm_reduce_add3b0_xor3b_wx125;
  wire multm_reduce_add3b0_xor3b_wx126;
  wire multm_reduce_add3b0_xor3b_wx127;
  wire multm_reduce_add3b0_xor3b_wx128;
  wire multm_reduce_add3b0_xor3b_wx129;
  wire multm_reduce_add3b0_xor3b_wx130;
  wire multm_reduce_add3b0_xor3b_wx131;
  wire multm_reduce_add3b0_xor3b_wx132;
  wire multm_reduce_add3b0_xor3b_wx133;
  wire multm_reduce_add3b0_xor3b_wx134;
  wire multm_reduce_add3b0_xor3b_wx135;
  wire multm_reduce_add3b0_xor3b_wx136;
  wire multm_reduce_add3b0_xor3b_wx137;
  wire multm_reduce_add3b0_xor3b_wx138;
  wire multm_reduce_add3b0_xor3b_wx139;
  wire multm_reduce_add3b0_xor3b_wx140;
  wire multm_reduce_add3b0_xor3b_wx141;
  wire multm_reduce_add3b0_xor3b_wx142;
  wire multm_reduce_add3b0_xor3b_wx143;
  wire multm_reduce_add3b0_xor3b_wx144;
  wire multm_reduce_add3b0_xor3b_wx145;
  wire multm_reduce_add3b0_xor3b_wx146;
  wire multm_reduce_add3b0_xor3b_wx147;
  wire multm_reduce_add3b0_xor3b_wx148;
  wire multm_reduce_add3b0_xor3b_wx149;
  wire multm_reduce_add3b0_xor3b_wx150;
  wire multm_reduce_add3b0_xor3b_wx151;
  wire multm_reduce_add3b0_xor3b_wx152;
  wire multm_reduce_add3b0_xor3b_wx153;
  wire multm_reduce_add3b0_xor3b_wx154;
  wire multm_reduce_add3b0_xor3b_wx155;
  wire multm_reduce_add3b0_xor3b_wx156;
  wire multm_reduce_add3b0_xor3b_wx157;
  wire multm_reduce_add3b0_xor3b_wx158;
  wire multm_reduce_add3b0_xor3b_wx159;
  wire multm_reduce_add3b0_xor3b_wx160;
  wire multm_reduce_add3b0_xor3b_wx161;
  wire multm_reduce_add3b0_xor3b_wx162;
  wire multm_reduce_add3b0_xor3b_wx163;
  wire multm_reduce_add3b0_xor3b_wx164;
  wire multm_reduce_add3b0_xor3b_wx165;
  wire multm_reduce_add3b0_xor3b_wx166;
  wire multm_reduce_add3b0_xor3b_wx167;
  wire multm_reduce_add3b0_xor3b_wx168;
  wire multm_reduce_add3b0_xor3b_wx169;
  wire multm_reduce_add3b0_xor3b_wx170;
  wire multm_reduce_add3b0_xor3b_wx171;
  wire multm_reduce_add3b0_xor3b_wx172;
  wire multm_reduce_add3b0_xor3b_wx173;
  wire multm_reduce_add3b0_xor3b_wx174;
  wire multm_reduce_add3b0_xor3b_wx175;
  wire multm_reduce_add3b0_xor3b_wx176;
  wire multm_reduce_add3b0_xor3b_wx177;
  wire multm_reduce_add3b0_xor3b_wx178;
  wire multm_reduce_add3b0_xor3b_wx179;
  wire multm_reduce_add3b0_xor3b_wx180;
  wire multm_reduce_add3b0_xor3b_wx181;
  wire multm_reduce_add3b0_xor3b_wx182;
  wire multm_reduce_add3b1_maj3b_or3b_wx0;
  wire multm_reduce_add3b1_maj3b_or3b_wx1;
  wire multm_reduce_add3b1_maj3b_or3b_wx2;
  wire multm_reduce_add3b1_maj3b_or3b_wx3;
  wire multm_reduce_add3b1_maj3b_or3b_wx4;
  wire multm_reduce_add3b1_maj3b_or3b_wx5;
  wire multm_reduce_add3b1_maj3b_or3b_wx6;
  wire multm_reduce_add3b1_maj3b_or3b_wx7;
  wire multm_reduce_add3b1_maj3b_or3b_wx8;
  wire multm_reduce_add3b1_maj3b_or3b_wx9;
  wire multm_reduce_add3b1_maj3b_or3b_wx10;
  wire multm_reduce_add3b1_maj3b_or3b_wx11;
  wire multm_reduce_add3b1_maj3b_or3b_wx12;
  wire multm_reduce_add3b1_maj3b_or3b_wx13;
  wire multm_reduce_add3b1_maj3b_or3b_wx14;
  wire multm_reduce_add3b1_maj3b_or3b_wx15;
  wire multm_reduce_add3b1_maj3b_or3b_wx16;
  wire multm_reduce_add3b1_maj3b_or3b_wx17;
  wire multm_reduce_add3b1_maj3b_or3b_wx18;
  wire multm_reduce_add3b1_maj3b_or3b_wx19;
  wire multm_reduce_add3b1_maj3b_or3b_wx20;
  wire multm_reduce_add3b1_maj3b_or3b_wx21;
  wire multm_reduce_add3b1_maj3b_or3b_wx22;
  wire multm_reduce_add3b1_maj3b_or3b_wx23;
  wire multm_reduce_add3b1_maj3b_or3b_wx24;
  wire multm_reduce_add3b1_maj3b_or3b_wx25;
  wire multm_reduce_add3b1_maj3b_or3b_wx26;
  wire multm_reduce_add3b1_maj3b_or3b_wx27;
  wire multm_reduce_add3b1_maj3b_or3b_wx28;
  wire multm_reduce_add3b1_maj3b_or3b_wx29;
  wire multm_reduce_add3b1_maj3b_or3b_wx30;
  wire multm_reduce_add3b1_maj3b_or3b_wx31;
  wire multm_reduce_add3b1_maj3b_or3b_wx32;
  wire multm_reduce_add3b1_maj3b_or3b_wx33;
  wire multm_reduce_add3b1_maj3b_or3b_wx34;
  wire multm_reduce_add3b1_maj3b_or3b_wx35;
  wire multm_reduce_add3b1_maj3b_or3b_wx36;
  wire multm_reduce_add3b1_maj3b_or3b_wx37;
  wire multm_reduce_add3b1_maj3b_or3b_wx38;
  wire multm_reduce_add3b1_maj3b_or3b_wx39;
  wire multm_reduce_add3b1_maj3b_or3b_wx40;
  wire multm_reduce_add3b1_maj3b_or3b_wx41;
  wire multm_reduce_add3b1_maj3b_or3b_wx42;
  wire multm_reduce_add3b1_maj3b_or3b_wx43;
  wire multm_reduce_add3b1_maj3b_or3b_wx44;
  wire multm_reduce_add3b1_maj3b_or3b_wx45;
  wire multm_reduce_add3b1_maj3b_or3b_wx46;
  wire multm_reduce_add3b1_maj3b_or3b_wx47;
  wire multm_reduce_add3b1_maj3b_or3b_wx48;
  wire multm_reduce_add3b1_maj3b_or3b_wx49;
  wire multm_reduce_add3b1_maj3b_or3b_wx50;
  wire multm_reduce_add3b1_maj3b_or3b_wx51;
  wire multm_reduce_add3b1_maj3b_or3b_wx52;
  wire multm_reduce_add3b1_maj3b_or3b_wx53;
  wire multm_reduce_add3b1_maj3b_or3b_wx54;
  wire multm_reduce_add3b1_maj3b_or3b_wx55;
  wire multm_reduce_add3b1_maj3b_or3b_wx56;
  wire multm_reduce_add3b1_maj3b_or3b_wx57;
  wire multm_reduce_add3b1_maj3b_or3b_wx58;
  wire multm_reduce_add3b1_maj3b_or3b_wx59;
  wire multm_reduce_add3b1_maj3b_or3b_wx60;
  wire multm_reduce_add3b1_maj3b_or3b_wx61;
  wire multm_reduce_add3b1_maj3b_or3b_wx62;
  wire multm_reduce_add3b1_maj3b_or3b_wx63;
  wire multm_reduce_add3b1_maj3b_or3b_wx64;
  wire multm_reduce_add3b1_maj3b_or3b_wx65;
  wire multm_reduce_add3b1_maj3b_or3b_wx66;
  wire multm_reduce_add3b1_maj3b_or3b_wx67;
  wire multm_reduce_add3b1_maj3b_or3b_wx68;
  wire multm_reduce_add3b1_maj3b_or3b_wx69;
  wire multm_reduce_add3b1_maj3b_or3b_wx70;
  wire multm_reduce_add3b1_maj3b_or3b_wx71;
  wire multm_reduce_add3b1_maj3b_or3b_wx72;
  wire multm_reduce_add3b1_maj3b_or3b_wx73;
  wire multm_reduce_add3b1_maj3b_or3b_wx74;
  wire multm_reduce_add3b1_maj3b_or3b_wx75;
  wire multm_reduce_add3b1_maj3b_or3b_wx76;
  wire multm_reduce_add3b1_maj3b_or3b_wx77;
  wire multm_reduce_add3b1_maj3b_or3b_wx78;
  wire multm_reduce_add3b1_maj3b_or3b_wx79;
  wire multm_reduce_add3b1_maj3b_or3b_wx80;
  wire multm_reduce_add3b1_maj3b_or3b_wx81;
  wire multm_reduce_add3b1_maj3b_or3b_wx82;
  wire multm_reduce_add3b1_maj3b_or3b_wx83;
  wire multm_reduce_add3b1_maj3b_or3b_wx84;
  wire multm_reduce_add3b1_maj3b_or3b_wx85;
  wire multm_reduce_add3b1_maj3b_or3b_wx86;
  wire multm_reduce_add3b1_maj3b_or3b_wx87;
  wire multm_reduce_add3b1_maj3b_or3b_wx88;
  wire multm_reduce_add3b1_maj3b_or3b_wx89;
  wire multm_reduce_add3b1_maj3b_or3b_wx90;
  wire multm_reduce_add3b1_maj3b_or3b_wx91;
  wire multm_reduce_add3b1_maj3b_or3b_wx92;
  wire multm_reduce_add3b1_maj3b_or3b_wx93;
  wire multm_reduce_add3b1_maj3b_or3b_wx94;
  wire multm_reduce_add3b1_maj3b_or3b_wx95;
  wire multm_reduce_add3b1_maj3b_or3b_wx96;
  wire multm_reduce_add3b1_maj3b_or3b_wx97;
  wire multm_reduce_add3b1_maj3b_or3b_wx98;
  wire multm_reduce_add3b1_maj3b_or3b_wx99;
  wire multm_reduce_add3b1_maj3b_or3b_wx100;
  wire multm_reduce_add3b1_maj3b_or3b_wx101;
  wire multm_reduce_add3b1_maj3b_or3b_wx102;
  wire multm_reduce_add3b1_maj3b_or3b_wx103;
  wire multm_reduce_add3b1_maj3b_or3b_wx104;
  wire multm_reduce_add3b1_maj3b_or3b_wx105;
  wire multm_reduce_add3b1_maj3b_or3b_wx106;
  wire multm_reduce_add3b1_maj3b_or3b_wx107;
  wire multm_reduce_add3b1_maj3b_or3b_wx108;
  wire multm_reduce_add3b1_maj3b_or3b_wx109;
  wire multm_reduce_add3b1_maj3b_or3b_wx110;
  wire multm_reduce_add3b1_maj3b_or3b_wx111;
  wire multm_reduce_add3b1_maj3b_or3b_wx112;
  wire multm_reduce_add3b1_maj3b_or3b_wx113;
  wire multm_reduce_add3b1_maj3b_or3b_wx114;
  wire multm_reduce_add3b1_maj3b_or3b_wx115;
  wire multm_reduce_add3b1_maj3b_or3b_wx116;
  wire multm_reduce_add3b1_maj3b_or3b_wx117;
  wire multm_reduce_add3b1_maj3b_or3b_wx118;
  wire multm_reduce_add3b1_maj3b_or3b_wx119;
  wire multm_reduce_add3b1_maj3b_or3b_wx120;
  wire multm_reduce_add3b1_maj3b_or3b_wx121;
  wire multm_reduce_add3b1_maj3b_or3b_wx122;
  wire multm_reduce_add3b1_maj3b_or3b_wx123;
  wire multm_reduce_add3b1_maj3b_or3b_wx124;
  wire multm_reduce_add3b1_maj3b_or3b_wx125;
  wire multm_reduce_add3b1_maj3b_or3b_wx126;
  wire multm_reduce_add3b1_maj3b_or3b_wx127;
  wire multm_reduce_add3b1_maj3b_or3b_wx128;
  wire multm_reduce_add3b1_maj3b_or3b_wx129;
  wire multm_reduce_add3b1_maj3b_or3b_wx130;
  wire multm_reduce_add3b1_maj3b_or3b_wx131;
  wire multm_reduce_add3b1_maj3b_or3b_wx132;
  wire multm_reduce_add3b1_maj3b_or3b_wx133;
  wire multm_reduce_add3b1_maj3b_or3b_wx134;
  wire multm_reduce_add3b1_maj3b_or3b_wx135;
  wire multm_reduce_add3b1_maj3b_or3b_wx136;
  wire multm_reduce_add3b1_maj3b_or3b_wx137;
  wire multm_reduce_add3b1_maj3b_or3b_wx138;
  wire multm_reduce_add3b1_maj3b_or3b_wx139;
  wire multm_reduce_add3b1_maj3b_or3b_wx140;
  wire multm_reduce_add3b1_maj3b_or3b_wx141;
  wire multm_reduce_add3b1_maj3b_or3b_wx142;
  wire multm_reduce_add3b1_maj3b_or3b_wx143;
  wire multm_reduce_add3b1_maj3b_or3b_wx144;
  wire multm_reduce_add3b1_maj3b_or3b_wx145;
  wire multm_reduce_add3b1_maj3b_or3b_wx146;
  wire multm_reduce_add3b1_maj3b_or3b_wx147;
  wire multm_reduce_add3b1_maj3b_or3b_wx148;
  wire multm_reduce_add3b1_maj3b_or3b_wx149;
  wire multm_reduce_add3b1_maj3b_or3b_wx150;
  wire multm_reduce_add3b1_maj3b_or3b_wx151;
  wire multm_reduce_add3b1_maj3b_or3b_wx152;
  wire multm_reduce_add3b1_maj3b_or3b_wx153;
  wire multm_reduce_add3b1_maj3b_or3b_wx154;
  wire multm_reduce_add3b1_maj3b_or3b_wx155;
  wire multm_reduce_add3b1_maj3b_or3b_wx156;
  wire multm_reduce_add3b1_maj3b_or3b_wx157;
  wire multm_reduce_add3b1_maj3b_or3b_wx158;
  wire multm_reduce_add3b1_maj3b_or3b_wx159;
  wire multm_reduce_add3b1_maj3b_or3b_wx160;
  wire multm_reduce_add3b1_maj3b_or3b_wx161;
  wire multm_reduce_add3b1_maj3b_or3b_wx162;
  wire multm_reduce_add3b1_maj3b_or3b_wx163;
  wire multm_reduce_add3b1_maj3b_or3b_wx164;
  wire multm_reduce_add3b1_maj3b_or3b_wx165;
  wire multm_reduce_add3b1_maj3b_or3b_wx166;
  wire multm_reduce_add3b1_maj3b_or3b_wx167;
  wire multm_reduce_add3b1_maj3b_or3b_wx168;
  wire multm_reduce_add3b1_maj3b_or3b_wx169;
  wire multm_reduce_add3b1_maj3b_or3b_wx170;
  wire multm_reduce_add3b1_maj3b_or3b_wx171;
  wire multm_reduce_add3b1_maj3b_or3b_wx172;
  wire multm_reduce_add3b1_maj3b_wx0;
  wire multm_reduce_add3b1_maj3b_wx1;
  wire multm_reduce_add3b1_maj3b_wx2;
  wire multm_reduce_add3b1_maj3b_wx3;
  wire multm_reduce_add3b1_maj3b_wx4;
  wire multm_reduce_add3b1_maj3b_wx5;
  wire multm_reduce_add3b1_maj3b_wx6;
  wire multm_reduce_add3b1_maj3b_wx7;
  wire multm_reduce_add3b1_maj3b_wx8;
  wire multm_reduce_add3b1_maj3b_wx9;
  wire multm_reduce_add3b1_maj3b_wx10;
  wire multm_reduce_add3b1_maj3b_wx11;
  wire multm_reduce_add3b1_maj3b_wx12;
  wire multm_reduce_add3b1_maj3b_wx13;
  wire multm_reduce_add3b1_maj3b_wx14;
  wire multm_reduce_add3b1_maj3b_wx15;
  wire multm_reduce_add3b1_maj3b_wx16;
  wire multm_reduce_add3b1_maj3b_wx17;
  wire multm_reduce_add3b1_maj3b_wx18;
  wire multm_reduce_add3b1_maj3b_wx19;
  wire multm_reduce_add3b1_maj3b_wx20;
  wire multm_reduce_add3b1_maj3b_wx21;
  wire multm_reduce_add3b1_maj3b_wx22;
  wire multm_reduce_add3b1_maj3b_wx23;
  wire multm_reduce_add3b1_maj3b_wx24;
  wire multm_reduce_add3b1_maj3b_wx25;
  wire multm_reduce_add3b1_maj3b_wx26;
  wire multm_reduce_add3b1_maj3b_wx27;
  wire multm_reduce_add3b1_maj3b_wx28;
  wire multm_reduce_add3b1_maj3b_wx29;
  wire multm_reduce_add3b1_maj3b_wx30;
  wire multm_reduce_add3b1_maj3b_wx31;
  wire multm_reduce_add3b1_maj3b_wx32;
  wire multm_reduce_add3b1_maj3b_wx33;
  wire multm_reduce_add3b1_maj3b_wx34;
  wire multm_reduce_add3b1_maj3b_wx35;
  wire multm_reduce_add3b1_maj3b_wx36;
  wire multm_reduce_add3b1_maj3b_wx37;
  wire multm_reduce_add3b1_maj3b_wx38;
  wire multm_reduce_add3b1_maj3b_wx39;
  wire multm_reduce_add3b1_maj3b_wx40;
  wire multm_reduce_add3b1_maj3b_wx41;
  wire multm_reduce_add3b1_maj3b_wx42;
  wire multm_reduce_add3b1_maj3b_wx43;
  wire multm_reduce_add3b1_maj3b_wx44;
  wire multm_reduce_add3b1_maj3b_wx45;
  wire multm_reduce_add3b1_maj3b_wx46;
  wire multm_reduce_add3b1_maj3b_wx47;
  wire multm_reduce_add3b1_maj3b_wx48;
  wire multm_reduce_add3b1_maj3b_wx49;
  wire multm_reduce_add3b1_maj3b_wx50;
  wire multm_reduce_add3b1_maj3b_wx51;
  wire multm_reduce_add3b1_maj3b_wx52;
  wire multm_reduce_add3b1_maj3b_wx53;
  wire multm_reduce_add3b1_maj3b_wx54;
  wire multm_reduce_add3b1_maj3b_wx55;
  wire multm_reduce_add3b1_maj3b_wx56;
  wire multm_reduce_add3b1_maj3b_wx57;
  wire multm_reduce_add3b1_maj3b_wx58;
  wire multm_reduce_add3b1_maj3b_wx59;
  wire multm_reduce_add3b1_maj3b_wx60;
  wire multm_reduce_add3b1_maj3b_wx61;
  wire multm_reduce_add3b1_maj3b_wx62;
  wire multm_reduce_add3b1_maj3b_wx63;
  wire multm_reduce_add3b1_maj3b_wx64;
  wire multm_reduce_add3b1_maj3b_wx65;
  wire multm_reduce_add3b1_maj3b_wx66;
  wire multm_reduce_add3b1_maj3b_wx67;
  wire multm_reduce_add3b1_maj3b_wx68;
  wire multm_reduce_add3b1_maj3b_wx69;
  wire multm_reduce_add3b1_maj3b_wx70;
  wire multm_reduce_add3b1_maj3b_wx71;
  wire multm_reduce_add3b1_maj3b_wx72;
  wire multm_reduce_add3b1_maj3b_wx73;
  wire multm_reduce_add3b1_maj3b_wx74;
  wire multm_reduce_add3b1_maj3b_wx75;
  wire multm_reduce_add3b1_maj3b_wx76;
  wire multm_reduce_add3b1_maj3b_wx77;
  wire multm_reduce_add3b1_maj3b_wx78;
  wire multm_reduce_add3b1_maj3b_wx79;
  wire multm_reduce_add3b1_maj3b_wx80;
  wire multm_reduce_add3b1_maj3b_wx81;
  wire multm_reduce_add3b1_maj3b_wx82;
  wire multm_reduce_add3b1_maj3b_wx83;
  wire multm_reduce_add3b1_maj3b_wx84;
  wire multm_reduce_add3b1_maj3b_wx85;
  wire multm_reduce_add3b1_maj3b_wx86;
  wire multm_reduce_add3b1_maj3b_wx87;
  wire multm_reduce_add3b1_maj3b_wx88;
  wire multm_reduce_add3b1_maj3b_wx89;
  wire multm_reduce_add3b1_maj3b_wx90;
  wire multm_reduce_add3b1_maj3b_wx91;
  wire multm_reduce_add3b1_maj3b_wx92;
  wire multm_reduce_add3b1_maj3b_wx93;
  wire multm_reduce_add3b1_maj3b_wx94;
  wire multm_reduce_add3b1_maj3b_wx95;
  wire multm_reduce_add3b1_maj3b_wx96;
  wire multm_reduce_add3b1_maj3b_wx97;
  wire multm_reduce_add3b1_maj3b_wx98;
  wire multm_reduce_add3b1_maj3b_wx99;
  wire multm_reduce_add3b1_maj3b_wx100;
  wire multm_reduce_add3b1_maj3b_wx101;
  wire multm_reduce_add3b1_maj3b_wx102;
  wire multm_reduce_add3b1_maj3b_wx103;
  wire multm_reduce_add3b1_maj3b_wx104;
  wire multm_reduce_add3b1_maj3b_wx105;
  wire multm_reduce_add3b1_maj3b_wx106;
  wire multm_reduce_add3b1_maj3b_wx107;
  wire multm_reduce_add3b1_maj3b_wx108;
  wire multm_reduce_add3b1_maj3b_wx109;
  wire multm_reduce_add3b1_maj3b_wx110;
  wire multm_reduce_add3b1_maj3b_wx111;
  wire multm_reduce_add3b1_maj3b_wx112;
  wire multm_reduce_add3b1_maj3b_wx113;
  wire multm_reduce_add3b1_maj3b_wx114;
  wire multm_reduce_add3b1_maj3b_wx115;
  wire multm_reduce_add3b1_maj3b_wx116;
  wire multm_reduce_add3b1_maj3b_wx117;
  wire multm_reduce_add3b1_maj3b_wx118;
  wire multm_reduce_add3b1_maj3b_wx119;
  wire multm_reduce_add3b1_maj3b_wx120;
  wire multm_reduce_add3b1_maj3b_wx121;
  wire multm_reduce_add3b1_maj3b_wx122;
  wire multm_reduce_add3b1_maj3b_wx123;
  wire multm_reduce_add3b1_maj3b_wx124;
  wire multm_reduce_add3b1_maj3b_wx125;
  wire multm_reduce_add3b1_maj3b_wx126;
  wire multm_reduce_add3b1_maj3b_wx127;
  wire multm_reduce_add3b1_maj3b_wx128;
  wire multm_reduce_add3b1_maj3b_wx129;
  wire multm_reduce_add3b1_maj3b_wx130;
  wire multm_reduce_add3b1_maj3b_wx131;
  wire multm_reduce_add3b1_maj3b_wx132;
  wire multm_reduce_add3b1_maj3b_wx133;
  wire multm_reduce_add3b1_maj3b_wx134;
  wire multm_reduce_add3b1_maj3b_wx135;
  wire multm_reduce_add3b1_maj3b_wx136;
  wire multm_reduce_add3b1_maj3b_wx137;
  wire multm_reduce_add3b1_maj3b_wx138;
  wire multm_reduce_add3b1_maj3b_wx139;
  wire multm_reduce_add3b1_maj3b_wx140;
  wire multm_reduce_add3b1_maj3b_wx141;
  wire multm_reduce_add3b1_maj3b_wx142;
  wire multm_reduce_add3b1_maj3b_wx143;
  wire multm_reduce_add3b1_maj3b_wx144;
  wire multm_reduce_add3b1_maj3b_wx145;
  wire multm_reduce_add3b1_maj3b_wx146;
  wire multm_reduce_add3b1_maj3b_wx147;
  wire multm_reduce_add3b1_maj3b_wx148;
  wire multm_reduce_add3b1_maj3b_wx149;
  wire multm_reduce_add3b1_maj3b_wx150;
  wire multm_reduce_add3b1_maj3b_wx151;
  wire multm_reduce_add3b1_maj3b_wx152;
  wire multm_reduce_add3b1_maj3b_wx153;
  wire multm_reduce_add3b1_maj3b_wx154;
  wire multm_reduce_add3b1_maj3b_wx155;
  wire multm_reduce_add3b1_maj3b_wx156;
  wire multm_reduce_add3b1_maj3b_wx157;
  wire multm_reduce_add3b1_maj3b_wx158;
  wire multm_reduce_add3b1_maj3b_wx159;
  wire multm_reduce_add3b1_maj3b_wx160;
  wire multm_reduce_add3b1_maj3b_wx161;
  wire multm_reduce_add3b1_maj3b_wx162;
  wire multm_reduce_add3b1_maj3b_wx163;
  wire multm_reduce_add3b1_maj3b_wx164;
  wire multm_reduce_add3b1_maj3b_wx165;
  wire multm_reduce_add3b1_maj3b_wx166;
  wire multm_reduce_add3b1_maj3b_wx167;
  wire multm_reduce_add3b1_maj3b_wx168;
  wire multm_reduce_add3b1_maj3b_wx169;
  wire multm_reduce_add3b1_maj3b_wx170;
  wire multm_reduce_add3b1_maj3b_wx171;
  wire multm_reduce_add3b1_maj3b_wx172;
  wire multm_reduce_add3b1_maj3b_wy0;
  wire multm_reduce_add3b1_maj3b_wy1;
  wire multm_reduce_add3b1_maj3b_wy2;
  wire multm_reduce_add3b1_maj3b_wy3;
  wire multm_reduce_add3b1_maj3b_wy4;
  wire multm_reduce_add3b1_maj3b_wy5;
  wire multm_reduce_add3b1_maj3b_wy6;
  wire multm_reduce_add3b1_maj3b_wy7;
  wire multm_reduce_add3b1_maj3b_wy8;
  wire multm_reduce_add3b1_maj3b_wy9;
  wire multm_reduce_add3b1_maj3b_wy10;
  wire multm_reduce_add3b1_maj3b_wy11;
  wire multm_reduce_add3b1_maj3b_wy12;
  wire multm_reduce_add3b1_maj3b_wy13;
  wire multm_reduce_add3b1_maj3b_wy14;
  wire multm_reduce_add3b1_maj3b_wy15;
  wire multm_reduce_add3b1_maj3b_wy16;
  wire multm_reduce_add3b1_maj3b_wy17;
  wire multm_reduce_add3b1_maj3b_wy18;
  wire multm_reduce_add3b1_maj3b_wy19;
  wire multm_reduce_add3b1_maj3b_wy20;
  wire multm_reduce_add3b1_maj3b_wy21;
  wire multm_reduce_add3b1_maj3b_wy22;
  wire multm_reduce_add3b1_maj3b_wy23;
  wire multm_reduce_add3b1_maj3b_wy24;
  wire multm_reduce_add3b1_maj3b_wy25;
  wire multm_reduce_add3b1_maj3b_wy26;
  wire multm_reduce_add3b1_maj3b_wy27;
  wire multm_reduce_add3b1_maj3b_wy28;
  wire multm_reduce_add3b1_maj3b_wy29;
  wire multm_reduce_add3b1_maj3b_wy30;
  wire multm_reduce_add3b1_maj3b_wy31;
  wire multm_reduce_add3b1_maj3b_wy32;
  wire multm_reduce_add3b1_maj3b_wy33;
  wire multm_reduce_add3b1_maj3b_wy34;
  wire multm_reduce_add3b1_maj3b_wy35;
  wire multm_reduce_add3b1_maj3b_wy36;
  wire multm_reduce_add3b1_maj3b_wy37;
  wire multm_reduce_add3b1_maj3b_wy38;
  wire multm_reduce_add3b1_maj3b_wy39;
  wire multm_reduce_add3b1_maj3b_wy40;
  wire multm_reduce_add3b1_maj3b_wy41;
  wire multm_reduce_add3b1_maj3b_wy42;
  wire multm_reduce_add3b1_maj3b_wy43;
  wire multm_reduce_add3b1_maj3b_wy44;
  wire multm_reduce_add3b1_maj3b_wy45;
  wire multm_reduce_add3b1_maj3b_wy46;
  wire multm_reduce_add3b1_maj3b_wy47;
  wire multm_reduce_add3b1_maj3b_wy48;
  wire multm_reduce_add3b1_maj3b_wy49;
  wire multm_reduce_add3b1_maj3b_wy50;
  wire multm_reduce_add3b1_maj3b_wy51;
  wire multm_reduce_add3b1_maj3b_wy52;
  wire multm_reduce_add3b1_maj3b_wy53;
  wire multm_reduce_add3b1_maj3b_wy54;
  wire multm_reduce_add3b1_maj3b_wy55;
  wire multm_reduce_add3b1_maj3b_wy56;
  wire multm_reduce_add3b1_maj3b_wy57;
  wire multm_reduce_add3b1_maj3b_wy58;
  wire multm_reduce_add3b1_maj3b_wy59;
  wire multm_reduce_add3b1_maj3b_wy60;
  wire multm_reduce_add3b1_maj3b_wy61;
  wire multm_reduce_add3b1_maj3b_wy62;
  wire multm_reduce_add3b1_maj3b_wy63;
  wire multm_reduce_add3b1_maj3b_wy64;
  wire multm_reduce_add3b1_maj3b_wy65;
  wire multm_reduce_add3b1_maj3b_wy66;
  wire multm_reduce_add3b1_maj3b_wy67;
  wire multm_reduce_add3b1_maj3b_wy68;
  wire multm_reduce_add3b1_maj3b_wy69;
  wire multm_reduce_add3b1_maj3b_wy70;
  wire multm_reduce_add3b1_maj3b_wy71;
  wire multm_reduce_add3b1_maj3b_wy72;
  wire multm_reduce_add3b1_maj3b_wy73;
  wire multm_reduce_add3b1_maj3b_wy74;
  wire multm_reduce_add3b1_maj3b_wy75;
  wire multm_reduce_add3b1_maj3b_wy76;
  wire multm_reduce_add3b1_maj3b_wy77;
  wire multm_reduce_add3b1_maj3b_wy78;
  wire multm_reduce_add3b1_maj3b_wy79;
  wire multm_reduce_add3b1_maj3b_wy80;
  wire multm_reduce_add3b1_maj3b_wy81;
  wire multm_reduce_add3b1_maj3b_wy82;
  wire multm_reduce_add3b1_maj3b_wy83;
  wire multm_reduce_add3b1_maj3b_wy84;
  wire multm_reduce_add3b1_maj3b_wy85;
  wire multm_reduce_add3b1_maj3b_wy86;
  wire multm_reduce_add3b1_maj3b_wy87;
  wire multm_reduce_add3b1_maj3b_wy88;
  wire multm_reduce_add3b1_maj3b_wy89;
  wire multm_reduce_add3b1_maj3b_wy90;
  wire multm_reduce_add3b1_maj3b_wy91;
  wire multm_reduce_add3b1_maj3b_wy92;
  wire multm_reduce_add3b1_maj3b_wy93;
  wire multm_reduce_add3b1_maj3b_wy94;
  wire multm_reduce_add3b1_maj3b_wy95;
  wire multm_reduce_add3b1_maj3b_wy96;
  wire multm_reduce_add3b1_maj3b_wy97;
  wire multm_reduce_add3b1_maj3b_wy98;
  wire multm_reduce_add3b1_maj3b_wy99;
  wire multm_reduce_add3b1_maj3b_wy100;
  wire multm_reduce_add3b1_maj3b_wy101;
  wire multm_reduce_add3b1_maj3b_wy102;
  wire multm_reduce_add3b1_maj3b_wy103;
  wire multm_reduce_add3b1_maj3b_wy104;
  wire multm_reduce_add3b1_maj3b_wy105;
  wire multm_reduce_add3b1_maj3b_wy106;
  wire multm_reduce_add3b1_maj3b_wy107;
  wire multm_reduce_add3b1_maj3b_wy108;
  wire multm_reduce_add3b1_maj3b_wy109;
  wire multm_reduce_add3b1_maj3b_wy110;
  wire multm_reduce_add3b1_maj3b_wy111;
  wire multm_reduce_add3b1_maj3b_wy112;
  wire multm_reduce_add3b1_maj3b_wy113;
  wire multm_reduce_add3b1_maj3b_wy114;
  wire multm_reduce_add3b1_maj3b_wy115;
  wire multm_reduce_add3b1_maj3b_wy116;
  wire multm_reduce_add3b1_maj3b_wy117;
  wire multm_reduce_add3b1_maj3b_wy118;
  wire multm_reduce_add3b1_maj3b_wy119;
  wire multm_reduce_add3b1_maj3b_wy120;
  wire multm_reduce_add3b1_maj3b_wy121;
  wire multm_reduce_add3b1_maj3b_wy122;
  wire multm_reduce_add3b1_maj3b_wy123;
  wire multm_reduce_add3b1_maj3b_wy124;
  wire multm_reduce_add3b1_maj3b_wy125;
  wire multm_reduce_add3b1_maj3b_wy126;
  wire multm_reduce_add3b1_maj3b_wy127;
  wire multm_reduce_add3b1_maj3b_wy128;
  wire multm_reduce_add3b1_maj3b_wy129;
  wire multm_reduce_add3b1_maj3b_wy130;
  wire multm_reduce_add3b1_maj3b_wy131;
  wire multm_reduce_add3b1_maj3b_wy132;
  wire multm_reduce_add3b1_maj3b_wy133;
  wire multm_reduce_add3b1_maj3b_wy134;
  wire multm_reduce_add3b1_maj3b_wy135;
  wire multm_reduce_add3b1_maj3b_wy136;
  wire multm_reduce_add3b1_maj3b_wy137;
  wire multm_reduce_add3b1_maj3b_wy138;
  wire multm_reduce_add3b1_maj3b_wy139;
  wire multm_reduce_add3b1_maj3b_wy140;
  wire multm_reduce_add3b1_maj3b_wy141;
  wire multm_reduce_add3b1_maj3b_wy142;
  wire multm_reduce_add3b1_maj3b_wy143;
  wire multm_reduce_add3b1_maj3b_wy144;
  wire multm_reduce_add3b1_maj3b_wy145;
  wire multm_reduce_add3b1_maj3b_wy146;
  wire multm_reduce_add3b1_maj3b_wy147;
  wire multm_reduce_add3b1_maj3b_wy148;
  wire multm_reduce_add3b1_maj3b_wy149;
  wire multm_reduce_add3b1_maj3b_wy150;
  wire multm_reduce_add3b1_maj3b_wy151;
  wire multm_reduce_add3b1_maj3b_wy152;
  wire multm_reduce_add3b1_maj3b_wy153;
  wire multm_reduce_add3b1_maj3b_wy154;
  wire multm_reduce_add3b1_maj3b_wy155;
  wire multm_reduce_add3b1_maj3b_wy156;
  wire multm_reduce_add3b1_maj3b_wy157;
  wire multm_reduce_add3b1_maj3b_wy158;
  wire multm_reduce_add3b1_maj3b_wy159;
  wire multm_reduce_add3b1_maj3b_wy160;
  wire multm_reduce_add3b1_maj3b_wy161;
  wire multm_reduce_add3b1_maj3b_wy162;
  wire multm_reduce_add3b1_maj3b_wy163;
  wire multm_reduce_add3b1_maj3b_wy164;
  wire multm_reduce_add3b1_maj3b_wy165;
  wire multm_reduce_add3b1_maj3b_wy166;
  wire multm_reduce_add3b1_maj3b_wy167;
  wire multm_reduce_add3b1_maj3b_wy168;
  wire multm_reduce_add3b1_maj3b_wy169;
  wire multm_reduce_add3b1_maj3b_wy170;
  wire multm_reduce_add3b1_maj3b_wy171;
  wire multm_reduce_add3b1_maj3b_wy172;
  wire multm_reduce_add3b1_maj3b_xy0;
  wire multm_reduce_add3b1_maj3b_xy1;
  wire multm_reduce_add3b1_maj3b_xy2;
  wire multm_reduce_add3b1_maj3b_xy3;
  wire multm_reduce_add3b1_maj3b_xy4;
  wire multm_reduce_add3b1_maj3b_xy5;
  wire multm_reduce_add3b1_maj3b_xy6;
  wire multm_reduce_add3b1_maj3b_xy7;
  wire multm_reduce_add3b1_maj3b_xy8;
  wire multm_reduce_add3b1_maj3b_xy9;
  wire multm_reduce_add3b1_maj3b_xy10;
  wire multm_reduce_add3b1_maj3b_xy11;
  wire multm_reduce_add3b1_maj3b_xy12;
  wire multm_reduce_add3b1_maj3b_xy13;
  wire multm_reduce_add3b1_maj3b_xy14;
  wire multm_reduce_add3b1_maj3b_xy15;
  wire multm_reduce_add3b1_maj3b_xy16;
  wire multm_reduce_add3b1_maj3b_xy17;
  wire multm_reduce_add3b1_maj3b_xy18;
  wire multm_reduce_add3b1_maj3b_xy19;
  wire multm_reduce_add3b1_maj3b_xy20;
  wire multm_reduce_add3b1_maj3b_xy21;
  wire multm_reduce_add3b1_maj3b_xy22;
  wire multm_reduce_add3b1_maj3b_xy23;
  wire multm_reduce_add3b1_maj3b_xy24;
  wire multm_reduce_add3b1_maj3b_xy25;
  wire multm_reduce_add3b1_maj3b_xy26;
  wire multm_reduce_add3b1_maj3b_xy27;
  wire multm_reduce_add3b1_maj3b_xy28;
  wire multm_reduce_add3b1_maj3b_xy29;
  wire multm_reduce_add3b1_maj3b_xy30;
  wire multm_reduce_add3b1_maj3b_xy31;
  wire multm_reduce_add3b1_maj3b_xy32;
  wire multm_reduce_add3b1_maj3b_xy33;
  wire multm_reduce_add3b1_maj3b_xy34;
  wire multm_reduce_add3b1_maj3b_xy35;
  wire multm_reduce_add3b1_maj3b_xy36;
  wire multm_reduce_add3b1_maj3b_xy37;
  wire multm_reduce_add3b1_maj3b_xy38;
  wire multm_reduce_add3b1_maj3b_xy39;
  wire multm_reduce_add3b1_maj3b_xy40;
  wire multm_reduce_add3b1_maj3b_xy41;
  wire multm_reduce_add3b1_maj3b_xy42;
  wire multm_reduce_add3b1_maj3b_xy43;
  wire multm_reduce_add3b1_maj3b_xy44;
  wire multm_reduce_add3b1_maj3b_xy45;
  wire multm_reduce_add3b1_maj3b_xy46;
  wire multm_reduce_add3b1_maj3b_xy47;
  wire multm_reduce_add3b1_maj3b_xy48;
  wire multm_reduce_add3b1_maj3b_xy49;
  wire multm_reduce_add3b1_maj3b_xy50;
  wire multm_reduce_add3b1_maj3b_xy51;
  wire multm_reduce_add3b1_maj3b_xy52;
  wire multm_reduce_add3b1_maj3b_xy53;
  wire multm_reduce_add3b1_maj3b_xy54;
  wire multm_reduce_add3b1_maj3b_xy55;
  wire multm_reduce_add3b1_maj3b_xy56;
  wire multm_reduce_add3b1_maj3b_xy57;
  wire multm_reduce_add3b1_maj3b_xy58;
  wire multm_reduce_add3b1_maj3b_xy59;
  wire multm_reduce_add3b1_maj3b_xy60;
  wire multm_reduce_add3b1_maj3b_xy61;
  wire multm_reduce_add3b1_maj3b_xy62;
  wire multm_reduce_add3b1_maj3b_xy63;
  wire multm_reduce_add3b1_maj3b_xy64;
  wire multm_reduce_add3b1_maj3b_xy65;
  wire multm_reduce_add3b1_maj3b_xy66;
  wire multm_reduce_add3b1_maj3b_xy67;
  wire multm_reduce_add3b1_maj3b_xy68;
  wire multm_reduce_add3b1_maj3b_xy69;
  wire multm_reduce_add3b1_maj3b_xy70;
  wire multm_reduce_add3b1_maj3b_xy71;
  wire multm_reduce_add3b1_maj3b_xy72;
  wire multm_reduce_add3b1_maj3b_xy73;
  wire multm_reduce_add3b1_maj3b_xy74;
  wire multm_reduce_add3b1_maj3b_xy75;
  wire multm_reduce_add3b1_maj3b_xy76;
  wire multm_reduce_add3b1_maj3b_xy77;
  wire multm_reduce_add3b1_maj3b_xy78;
  wire multm_reduce_add3b1_maj3b_xy79;
  wire multm_reduce_add3b1_maj3b_xy80;
  wire multm_reduce_add3b1_maj3b_xy81;
  wire multm_reduce_add3b1_maj3b_xy82;
  wire multm_reduce_add3b1_maj3b_xy83;
  wire multm_reduce_add3b1_maj3b_xy84;
  wire multm_reduce_add3b1_maj3b_xy85;
  wire multm_reduce_add3b1_maj3b_xy86;
  wire multm_reduce_add3b1_maj3b_xy87;
  wire multm_reduce_add3b1_maj3b_xy88;
  wire multm_reduce_add3b1_maj3b_xy89;
  wire multm_reduce_add3b1_maj3b_xy90;
  wire multm_reduce_add3b1_maj3b_xy91;
  wire multm_reduce_add3b1_maj3b_xy92;
  wire multm_reduce_add3b1_maj3b_xy93;
  wire multm_reduce_add3b1_maj3b_xy94;
  wire multm_reduce_add3b1_maj3b_xy95;
  wire multm_reduce_add3b1_maj3b_xy96;
  wire multm_reduce_add3b1_maj3b_xy97;
  wire multm_reduce_add3b1_maj3b_xy98;
  wire multm_reduce_add3b1_maj3b_xy99;
  wire multm_reduce_add3b1_maj3b_xy100;
  wire multm_reduce_add3b1_maj3b_xy101;
  wire multm_reduce_add3b1_maj3b_xy102;
  wire multm_reduce_add3b1_maj3b_xy103;
  wire multm_reduce_add3b1_maj3b_xy104;
  wire multm_reduce_add3b1_maj3b_xy105;
  wire multm_reduce_add3b1_maj3b_xy106;
  wire multm_reduce_add3b1_maj3b_xy107;
  wire multm_reduce_add3b1_maj3b_xy108;
  wire multm_reduce_add3b1_maj3b_xy109;
  wire multm_reduce_add3b1_maj3b_xy110;
  wire multm_reduce_add3b1_maj3b_xy111;
  wire multm_reduce_add3b1_maj3b_xy112;
  wire multm_reduce_add3b1_maj3b_xy113;
  wire multm_reduce_add3b1_maj3b_xy114;
  wire multm_reduce_add3b1_maj3b_xy115;
  wire multm_reduce_add3b1_maj3b_xy116;
  wire multm_reduce_add3b1_maj3b_xy117;
  wire multm_reduce_add3b1_maj3b_xy118;
  wire multm_reduce_add3b1_maj3b_xy119;
  wire multm_reduce_add3b1_maj3b_xy120;
  wire multm_reduce_add3b1_maj3b_xy121;
  wire multm_reduce_add3b1_maj3b_xy122;
  wire multm_reduce_add3b1_maj3b_xy123;
  wire multm_reduce_add3b1_maj3b_xy124;
  wire multm_reduce_add3b1_maj3b_xy125;
  wire multm_reduce_add3b1_maj3b_xy126;
  wire multm_reduce_add3b1_maj3b_xy127;
  wire multm_reduce_add3b1_maj3b_xy128;
  wire multm_reduce_add3b1_maj3b_xy129;
  wire multm_reduce_add3b1_maj3b_xy130;
  wire multm_reduce_add3b1_maj3b_xy131;
  wire multm_reduce_add3b1_maj3b_xy132;
  wire multm_reduce_add3b1_maj3b_xy133;
  wire multm_reduce_add3b1_maj3b_xy134;
  wire multm_reduce_add3b1_maj3b_xy135;
  wire multm_reduce_add3b1_maj3b_xy136;
  wire multm_reduce_add3b1_maj3b_xy137;
  wire multm_reduce_add3b1_maj3b_xy138;
  wire multm_reduce_add3b1_maj3b_xy139;
  wire multm_reduce_add3b1_maj3b_xy140;
  wire multm_reduce_add3b1_maj3b_xy141;
  wire multm_reduce_add3b1_maj3b_xy142;
  wire multm_reduce_add3b1_maj3b_xy143;
  wire multm_reduce_add3b1_maj3b_xy144;
  wire multm_reduce_add3b1_maj3b_xy145;
  wire multm_reduce_add3b1_maj3b_xy146;
  wire multm_reduce_add3b1_maj3b_xy147;
  wire multm_reduce_add3b1_maj3b_xy148;
  wire multm_reduce_add3b1_maj3b_xy149;
  wire multm_reduce_add3b1_maj3b_xy150;
  wire multm_reduce_add3b1_maj3b_xy151;
  wire multm_reduce_add3b1_maj3b_xy152;
  wire multm_reduce_add3b1_maj3b_xy153;
  wire multm_reduce_add3b1_maj3b_xy154;
  wire multm_reduce_add3b1_maj3b_xy155;
  wire multm_reduce_add3b1_maj3b_xy156;
  wire multm_reduce_add3b1_maj3b_xy157;
  wire multm_reduce_add3b1_maj3b_xy158;
  wire multm_reduce_add3b1_maj3b_xy159;
  wire multm_reduce_add3b1_maj3b_xy160;
  wire multm_reduce_add3b1_maj3b_xy161;
  wire multm_reduce_add3b1_maj3b_xy162;
  wire multm_reduce_add3b1_maj3b_xy163;
  wire multm_reduce_add3b1_maj3b_xy164;
  wire multm_reduce_add3b1_maj3b_xy165;
  wire multm_reduce_add3b1_maj3b_xy166;
  wire multm_reduce_add3b1_maj3b_xy167;
  wire multm_reduce_add3b1_maj3b_xy168;
  wire multm_reduce_add3b1_maj3b_xy169;
  wire multm_reduce_add3b1_maj3b_xy170;
  wire multm_reduce_add3b1_maj3b_xy171;
  wire multm_reduce_add3b1_maj3b_xy172;
  wire multm_reduce_add3b1_xor3b_wx0;
  wire multm_reduce_add3b1_xor3b_wx1;
  wire multm_reduce_add3b1_xor3b_wx2;
  wire multm_reduce_add3b1_xor3b_wx3;
  wire multm_reduce_add3b1_xor3b_wx4;
  wire multm_reduce_add3b1_xor3b_wx5;
  wire multm_reduce_add3b1_xor3b_wx6;
  wire multm_reduce_add3b1_xor3b_wx7;
  wire multm_reduce_add3b1_xor3b_wx8;
  wire multm_reduce_add3b1_xor3b_wx9;
  wire multm_reduce_add3b1_xor3b_wx10;
  wire multm_reduce_add3b1_xor3b_wx11;
  wire multm_reduce_add3b1_xor3b_wx12;
  wire multm_reduce_add3b1_xor3b_wx13;
  wire multm_reduce_add3b1_xor3b_wx14;
  wire multm_reduce_add3b1_xor3b_wx15;
  wire multm_reduce_add3b1_xor3b_wx16;
  wire multm_reduce_add3b1_xor3b_wx17;
  wire multm_reduce_add3b1_xor3b_wx18;
  wire multm_reduce_add3b1_xor3b_wx19;
  wire multm_reduce_add3b1_xor3b_wx20;
  wire multm_reduce_add3b1_xor3b_wx21;
  wire multm_reduce_add3b1_xor3b_wx22;
  wire multm_reduce_add3b1_xor3b_wx23;
  wire multm_reduce_add3b1_xor3b_wx24;
  wire multm_reduce_add3b1_xor3b_wx25;
  wire multm_reduce_add3b1_xor3b_wx26;
  wire multm_reduce_add3b1_xor3b_wx27;
  wire multm_reduce_add3b1_xor3b_wx28;
  wire multm_reduce_add3b1_xor3b_wx29;
  wire multm_reduce_add3b1_xor3b_wx30;
  wire multm_reduce_add3b1_xor3b_wx31;
  wire multm_reduce_add3b1_xor3b_wx32;
  wire multm_reduce_add3b1_xor3b_wx33;
  wire multm_reduce_add3b1_xor3b_wx34;
  wire multm_reduce_add3b1_xor3b_wx35;
  wire multm_reduce_add3b1_xor3b_wx36;
  wire multm_reduce_add3b1_xor3b_wx37;
  wire multm_reduce_add3b1_xor3b_wx38;
  wire multm_reduce_add3b1_xor3b_wx39;
  wire multm_reduce_add3b1_xor3b_wx40;
  wire multm_reduce_add3b1_xor3b_wx41;
  wire multm_reduce_add3b1_xor3b_wx42;
  wire multm_reduce_add3b1_xor3b_wx43;
  wire multm_reduce_add3b1_xor3b_wx44;
  wire multm_reduce_add3b1_xor3b_wx45;
  wire multm_reduce_add3b1_xor3b_wx46;
  wire multm_reduce_add3b1_xor3b_wx47;
  wire multm_reduce_add3b1_xor3b_wx48;
  wire multm_reduce_add3b1_xor3b_wx49;
  wire multm_reduce_add3b1_xor3b_wx50;
  wire multm_reduce_add3b1_xor3b_wx51;
  wire multm_reduce_add3b1_xor3b_wx52;
  wire multm_reduce_add3b1_xor3b_wx53;
  wire multm_reduce_add3b1_xor3b_wx54;
  wire multm_reduce_add3b1_xor3b_wx55;
  wire multm_reduce_add3b1_xor3b_wx56;
  wire multm_reduce_add3b1_xor3b_wx57;
  wire multm_reduce_add3b1_xor3b_wx58;
  wire multm_reduce_add3b1_xor3b_wx59;
  wire multm_reduce_add3b1_xor3b_wx60;
  wire multm_reduce_add3b1_xor3b_wx61;
  wire multm_reduce_add3b1_xor3b_wx62;
  wire multm_reduce_add3b1_xor3b_wx63;
  wire multm_reduce_add3b1_xor3b_wx64;
  wire multm_reduce_add3b1_xor3b_wx65;
  wire multm_reduce_add3b1_xor3b_wx66;
  wire multm_reduce_add3b1_xor3b_wx67;
  wire multm_reduce_add3b1_xor3b_wx68;
  wire multm_reduce_add3b1_xor3b_wx69;
  wire multm_reduce_add3b1_xor3b_wx70;
  wire multm_reduce_add3b1_xor3b_wx71;
  wire multm_reduce_add3b1_xor3b_wx72;
  wire multm_reduce_add3b1_xor3b_wx73;
  wire multm_reduce_add3b1_xor3b_wx74;
  wire multm_reduce_add3b1_xor3b_wx75;
  wire multm_reduce_add3b1_xor3b_wx76;
  wire multm_reduce_add3b1_xor3b_wx77;
  wire multm_reduce_add3b1_xor3b_wx78;
  wire multm_reduce_add3b1_xor3b_wx79;
  wire multm_reduce_add3b1_xor3b_wx80;
  wire multm_reduce_add3b1_xor3b_wx81;
  wire multm_reduce_add3b1_xor3b_wx82;
  wire multm_reduce_add3b1_xor3b_wx83;
  wire multm_reduce_add3b1_xor3b_wx84;
  wire multm_reduce_add3b1_xor3b_wx85;
  wire multm_reduce_add3b1_xor3b_wx86;
  wire multm_reduce_add3b1_xor3b_wx87;
  wire multm_reduce_add3b1_xor3b_wx88;
  wire multm_reduce_add3b1_xor3b_wx89;
  wire multm_reduce_add3b1_xor3b_wx90;
  wire multm_reduce_add3b1_xor3b_wx91;
  wire multm_reduce_add3b1_xor3b_wx92;
  wire multm_reduce_add3b1_xor3b_wx93;
  wire multm_reduce_add3b1_xor3b_wx94;
  wire multm_reduce_add3b1_xor3b_wx95;
  wire multm_reduce_add3b1_xor3b_wx96;
  wire multm_reduce_add3b1_xor3b_wx97;
  wire multm_reduce_add3b1_xor3b_wx98;
  wire multm_reduce_add3b1_xor3b_wx99;
  wire multm_reduce_add3b1_xor3b_wx100;
  wire multm_reduce_add3b1_xor3b_wx101;
  wire multm_reduce_add3b1_xor3b_wx102;
  wire multm_reduce_add3b1_xor3b_wx103;
  wire multm_reduce_add3b1_xor3b_wx104;
  wire multm_reduce_add3b1_xor3b_wx105;
  wire multm_reduce_add3b1_xor3b_wx106;
  wire multm_reduce_add3b1_xor3b_wx107;
  wire multm_reduce_add3b1_xor3b_wx108;
  wire multm_reduce_add3b1_xor3b_wx109;
  wire multm_reduce_add3b1_xor3b_wx110;
  wire multm_reduce_add3b1_xor3b_wx111;
  wire multm_reduce_add3b1_xor3b_wx112;
  wire multm_reduce_add3b1_xor3b_wx113;
  wire multm_reduce_add3b1_xor3b_wx114;
  wire multm_reduce_add3b1_xor3b_wx115;
  wire multm_reduce_add3b1_xor3b_wx116;
  wire multm_reduce_add3b1_xor3b_wx117;
  wire multm_reduce_add3b1_xor3b_wx118;
  wire multm_reduce_add3b1_xor3b_wx119;
  wire multm_reduce_add3b1_xor3b_wx120;
  wire multm_reduce_add3b1_xor3b_wx121;
  wire multm_reduce_add3b1_xor3b_wx122;
  wire multm_reduce_add3b1_xor3b_wx123;
  wire multm_reduce_add3b1_xor3b_wx124;
  wire multm_reduce_add3b1_xor3b_wx125;
  wire multm_reduce_add3b1_xor3b_wx126;
  wire multm_reduce_add3b1_xor3b_wx127;
  wire multm_reduce_add3b1_xor3b_wx128;
  wire multm_reduce_add3b1_xor3b_wx129;
  wire multm_reduce_add3b1_xor3b_wx130;
  wire multm_reduce_add3b1_xor3b_wx131;
  wire multm_reduce_add3b1_xor3b_wx132;
  wire multm_reduce_add3b1_xor3b_wx133;
  wire multm_reduce_add3b1_xor3b_wx134;
  wire multm_reduce_add3b1_xor3b_wx135;
  wire multm_reduce_add3b1_xor3b_wx136;
  wire multm_reduce_add3b1_xor3b_wx137;
  wire multm_reduce_add3b1_xor3b_wx138;
  wire multm_reduce_add3b1_xor3b_wx139;
  wire multm_reduce_add3b1_xor3b_wx140;
  wire multm_reduce_add3b1_xor3b_wx141;
  wire multm_reduce_add3b1_xor3b_wx142;
  wire multm_reduce_add3b1_xor3b_wx143;
  wire multm_reduce_add3b1_xor3b_wx144;
  wire multm_reduce_add3b1_xor3b_wx145;
  wire multm_reduce_add3b1_xor3b_wx146;
  wire multm_reduce_add3b1_xor3b_wx147;
  wire multm_reduce_add3b1_xor3b_wx148;
  wire multm_reduce_add3b1_xor3b_wx149;
  wire multm_reduce_add3b1_xor3b_wx150;
  wire multm_reduce_add3b1_xor3b_wx151;
  wire multm_reduce_add3b1_xor3b_wx152;
  wire multm_reduce_add3b1_xor3b_wx153;
  wire multm_reduce_add3b1_xor3b_wx154;
  wire multm_reduce_add3b1_xor3b_wx155;
  wire multm_reduce_add3b1_xor3b_wx156;
  wire multm_reduce_add3b1_xor3b_wx157;
  wire multm_reduce_add3b1_xor3b_wx158;
  wire multm_reduce_add3b1_xor3b_wx159;
  wire multm_reduce_add3b1_xor3b_wx160;
  wire multm_reduce_add3b1_xor3b_wx161;
  wire multm_reduce_add3b1_xor3b_wx162;
  wire multm_reduce_add3b1_xor3b_wx163;
  wire multm_reduce_add3b1_xor3b_wx164;
  wire multm_reduce_add3b1_xor3b_wx165;
  wire multm_reduce_add3b1_xor3b_wx166;
  wire multm_reduce_add3b1_xor3b_wx167;
  wire multm_reduce_add3b1_xor3b_wx168;
  wire multm_reduce_add3b1_xor3b_wx169;
  wire multm_reduce_add3b1_xor3b_wx170;
  wire multm_reduce_add3b1_xor3b_wx171;
  wire multm_reduce_add3b1_xor3b_wx172;
  wire multm_reduce_mc10;
  wire multm_reduce_mc11;
  wire multm_reduce_mc12;
  wire multm_reduce_mc13;
  wire multm_reduce_mc14;
  wire multm_reduce_mc15;
  wire multm_reduce_mc16;
  wire multm_reduce_mc17;
  wire multm_reduce_mc18;
  wire multm_reduce_mc19;
  wire multm_reduce_mc20;
  wire multm_reduce_mc21;
  wire multm_reduce_mc22;
  wire multm_reduce_mc23;
  wire multm_reduce_mc24;
  wire multm_reduce_mc25;
  wire multm_reduce_mc26;
  wire multm_reduce_mc27;
  wire multm_reduce_mc28;
  wire multm_reduce_mc29;
  wire multm_reduce_mc30;
  wire multm_reduce_mc31;
  wire multm_reduce_mc32;
  wire multm_reduce_mc33;
  wire multm_reduce_mc34;
  wire multm_reduce_mc35;
  wire multm_reduce_mc36;
  wire multm_reduce_mc37;
  wire multm_reduce_mc38;
  wire multm_reduce_mc39;
  wire multm_reduce_mc40;
  wire multm_reduce_mc41;
  wire multm_reduce_mc42;
  wire multm_reduce_mc43;
  wire multm_reduce_mc44;
  wire multm_reduce_mc45;
  wire multm_reduce_mc46;
  wire multm_reduce_mc47;
  wire multm_reduce_mc48;
  wire multm_reduce_mc49;
  wire multm_reduce_mc50;
  wire multm_reduce_mc51;
  wire multm_reduce_mc52;
  wire multm_reduce_mc53;
  wire multm_reduce_mc54;
  wire multm_reduce_mc55;
  wire multm_reduce_mc56;
  wire multm_reduce_mc57;
  wire multm_reduce_mc58;
  wire multm_reduce_mc59;
  wire multm_reduce_mc60;
  wire multm_reduce_mc61;
  wire multm_reduce_mc62;
  wire multm_reduce_mc63;
  wire multm_reduce_mc64;
  wire multm_reduce_mc65;
  wire multm_reduce_mc66;
  wire multm_reduce_mc67;
  wire multm_reduce_mc68;
  wire multm_reduce_mc69;
  wire multm_reduce_mc70;
  wire multm_reduce_mc71;
  wire multm_reduce_mc72;
  wire multm_reduce_mc73;
  wire multm_reduce_mc74;
  wire multm_reduce_mc75;
  wire multm_reduce_mc76;
  wire multm_reduce_mc77;
  wire multm_reduce_mc78;
  wire multm_reduce_mc79;
  wire multm_reduce_mc80;
  wire multm_reduce_mc81;
  wire multm_reduce_mc82;
  wire multm_reduce_mc83;
  wire multm_reduce_mc84;
  wire multm_reduce_mc85;
  wire multm_reduce_mc86;
  wire multm_reduce_mc87;
  wire multm_reduce_mc88;
  wire multm_reduce_mc89;
  wire multm_reduce_mc90;
  wire multm_reduce_mc91;
  wire multm_reduce_mc92;
  wire multm_reduce_mc93;
  wire multm_reduce_mc94;
  wire multm_reduce_mc95;
  wire multm_reduce_mc96;
  wire multm_reduce_mc97;
  wire multm_reduce_mc98;
  wire multm_reduce_mc99;
  wire multm_reduce_mc100;
  wire multm_reduce_mc101;
  wire multm_reduce_mc102;
  wire multm_reduce_mc103;
  wire multm_reduce_mc104;
  wire multm_reduce_mc105;
  wire multm_reduce_mc106;
  wire multm_reduce_mc107;
  wire multm_reduce_mc108;
  wire multm_reduce_mc109;
  wire multm_reduce_mc110;
  wire multm_reduce_mc111;
  wire multm_reduce_mc112;
  wire multm_reduce_mc113;
  wire multm_reduce_mc114;
  wire multm_reduce_mc115;
  wire multm_reduce_mc116;
  wire multm_reduce_mc117;
  wire multm_reduce_mc118;
  wire multm_reduce_mc119;
  wire multm_reduce_mc120;
  wire multm_reduce_mc121;
  wire multm_reduce_mc122;
  wire multm_reduce_mc123;
  wire multm_reduce_mc124;
  wire multm_reduce_mc125;
  wire multm_reduce_mc126;
  wire multm_reduce_mc127;
  wire multm_reduce_mc128;
  wire multm_reduce_mc129;
  wire multm_reduce_mc130;
  wire multm_reduce_mc131;
  wire multm_reduce_mc132;
  wire multm_reduce_mc133;
  wire multm_reduce_mc134;
  wire multm_reduce_mc135;
  wire multm_reduce_mc136;
  wire multm_reduce_mc137;
  wire multm_reduce_mc138;
  wire multm_reduce_mc139;
  wire multm_reduce_mc140;
  wire multm_reduce_mc141;
  wire multm_reduce_mc142;
  wire multm_reduce_mc143;
  wire multm_reduce_mc144;
  wire multm_reduce_mc145;
  wire multm_reduce_mc146;
  wire multm_reduce_mc147;
  wire multm_reduce_mc148;
  wire multm_reduce_mc149;
  wire multm_reduce_mc150;
  wire multm_reduce_mc151;
  wire multm_reduce_mc152;
  wire multm_reduce_mc153;
  wire multm_reduce_mc154;
  wire multm_reduce_mc155;
  wire multm_reduce_mc156;
  wire multm_reduce_mc157;
  wire multm_reduce_mc158;
  wire multm_reduce_mc159;
  wire multm_reduce_mc160;
  wire multm_reduce_mc161;
  wire multm_reduce_mc162;
  wire multm_reduce_mc163;
  wire multm_reduce_mc164;
  wire multm_reduce_mc165;
  wire multm_reduce_mc166;
  wire multm_reduce_mc167;
  wire multm_reduce_mc168;
  wire multm_reduce_mc169;
  wire multm_reduce_mc170;
  wire multm_reduce_mc171;
  wire multm_reduce_mc172;
  wire multm_reduce_mc173;
  wire multm_reduce_mc174;
  wire multm_reduce_mc175;
  wire multm_reduce_mc176;
  wire multm_reduce_mc177;
  wire multm_reduce_mc178;
  wire multm_reduce_mc179;
  wire multm_reduce_mc180;
  wire multm_reduce_mc181;
  wire multm_reduce_mc182;
  wire multm_reduce_mc183;
  wire multm_reduce_ms11;
  wire multm_reduce_ms12;
  wire multm_reduce_ms13;
  wire multm_reduce_ms14;
  wire multm_reduce_ms15;
  wire multm_reduce_ms16;
  wire multm_reduce_ms17;
  wire multm_reduce_ms18;
  wire multm_reduce_ms19;
  wire multm_reduce_ms20;
  wire multm_reduce_ms21;
  wire multm_reduce_ms22;
  wire multm_reduce_ms23;
  wire multm_reduce_ms24;
  wire multm_reduce_ms25;
  wire multm_reduce_ms26;
  wire multm_reduce_ms27;
  wire multm_reduce_ms28;
  wire multm_reduce_ms29;
  wire multm_reduce_ms30;
  wire multm_reduce_ms31;
  wire multm_reduce_ms32;
  wire multm_reduce_ms33;
  wire multm_reduce_ms34;
  wire multm_reduce_ms35;
  wire multm_reduce_ms36;
  wire multm_reduce_ms37;
  wire multm_reduce_ms38;
  wire multm_reduce_ms39;
  wire multm_reduce_ms40;
  wire multm_reduce_ms41;
  wire multm_reduce_ms42;
  wire multm_reduce_ms43;
  wire multm_reduce_ms44;
  wire multm_reduce_ms45;
  wire multm_reduce_ms46;
  wire multm_reduce_ms47;
  wire multm_reduce_ms48;
  wire multm_reduce_ms49;
  wire multm_reduce_ms50;
  wire multm_reduce_ms51;
  wire multm_reduce_ms52;
  wire multm_reduce_ms53;
  wire multm_reduce_ms54;
  wire multm_reduce_ms55;
  wire multm_reduce_ms56;
  wire multm_reduce_ms57;
  wire multm_reduce_ms58;
  wire multm_reduce_ms59;
  wire multm_reduce_ms60;
  wire multm_reduce_ms61;
  wire multm_reduce_ms62;
  wire multm_reduce_ms63;
  wire multm_reduce_ms64;
  wire multm_reduce_ms65;
  wire multm_reduce_ms66;
  wire multm_reduce_ms67;
  wire multm_reduce_ms68;
  wire multm_reduce_ms69;
  wire multm_reduce_ms70;
  wire multm_reduce_ms71;
  wire multm_reduce_ms72;
  wire multm_reduce_ms73;
  wire multm_reduce_ms74;
  wire multm_reduce_ms75;
  wire multm_reduce_ms76;
  wire multm_reduce_ms77;
  wire multm_reduce_ms78;
  wire multm_reduce_ms79;
  wire multm_reduce_ms80;
  wire multm_reduce_ms81;
  wire multm_reduce_ms82;
  wire multm_reduce_ms83;
  wire multm_reduce_ms84;
  wire multm_reduce_ms85;
  wire multm_reduce_ms86;
  wire multm_reduce_ms87;
  wire multm_reduce_ms88;
  wire multm_reduce_ms89;
  wire multm_reduce_ms90;
  wire multm_reduce_ms91;
  wire multm_reduce_ms92;
  wire multm_reduce_ms93;
  wire multm_reduce_ms94;
  wire multm_reduce_ms95;
  wire multm_reduce_ms96;
  wire multm_reduce_ms97;
  wire multm_reduce_ms98;
  wire multm_reduce_ms99;
  wire multm_reduce_ms100;
  wire multm_reduce_ms101;
  wire multm_reduce_ms102;
  wire multm_reduce_ms103;
  wire multm_reduce_ms104;
  wire multm_reduce_ms105;
  wire multm_reduce_ms106;
  wire multm_reduce_ms107;
  wire multm_reduce_ms108;
  wire multm_reduce_ms109;
  wire multm_reduce_ms110;
  wire multm_reduce_ms111;
  wire multm_reduce_ms112;
  wire multm_reduce_ms113;
  wire multm_reduce_ms114;
  wire multm_reduce_ms115;
  wire multm_reduce_ms116;
  wire multm_reduce_ms117;
  wire multm_reduce_ms118;
  wire multm_reduce_ms119;
  wire multm_reduce_ms120;
  wire multm_reduce_ms121;
  wire multm_reduce_ms122;
  wire multm_reduce_ms123;
  wire multm_reduce_ms124;
  wire multm_reduce_ms125;
  wire multm_reduce_ms126;
  wire multm_reduce_ms127;
  wire multm_reduce_ms128;
  wire multm_reduce_ms129;
  wire multm_reduce_ms130;
  wire multm_reduce_ms131;
  wire multm_reduce_ms132;
  wire multm_reduce_ms133;
  wire multm_reduce_ms134;
  wire multm_reduce_ms135;
  wire multm_reduce_ms136;
  wire multm_reduce_ms137;
  wire multm_reduce_ms138;
  wire multm_reduce_ms139;
  wire multm_reduce_ms140;
  wire multm_reduce_ms141;
  wire multm_reduce_ms142;
  wire multm_reduce_ms143;
  wire multm_reduce_ms144;
  wire multm_reduce_ms145;
  wire multm_reduce_ms146;
  wire multm_reduce_ms147;
  wire multm_reduce_ms148;
  wire multm_reduce_ms149;
  wire multm_reduce_ms150;
  wire multm_reduce_ms151;
  wire multm_reduce_ms152;
  wire multm_reduce_ms153;
  wire multm_reduce_ms154;
  wire multm_reduce_ms155;
  wire multm_reduce_ms156;
  wire multm_reduce_ms157;
  wire multm_reduce_ms158;
  wire multm_reduce_ms159;
  wire multm_reduce_ms160;
  wire multm_reduce_ms161;
  wire multm_reduce_ms162;
  wire multm_reduce_ms163;
  wire multm_reduce_ms164;
  wire multm_reduce_ms165;
  wire multm_reduce_ms166;
  wire multm_reduce_ms167;
  wire multm_reduce_ms168;
  wire multm_reduce_ms169;
  wire multm_reduce_ms170;
  wire multm_reduce_ms171;
  wire multm_reduce_ms172;
  wire multm_reduce_ms173;
  wire multm_reduce_ms174;
  wire multm_reduce_ms175;
  wire multm_reduce_ms176;
  wire multm_reduce_ms177;
  wire multm_reduce_ms178;
  wire multm_reduce_ms179;
  wire multm_reduce_ms180;
  wire multm_reduce_ms181;
  wire multm_reduce_ms182;
  wire multm_reduce_ms183;
  wire multm_reduce_mulb0_add3_maj3_or3_wx;
  wire multm_reduce_mulb0_add3_maj3_wx;
  wire multm_reduce_mulb0_add3_maj3_wy;
  wire multm_reduce_mulb0_add3_maj3_xy;
  wire multm_reduce_mulb0_add3_xor3_wx;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx2;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx4;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx8;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx9;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx12;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx15;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx16;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx17;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx18;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx19;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx20;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx25;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx26;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx27;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx29;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx30;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx33;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx37;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx40;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx42;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx44;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx45;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx46;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx48;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx50;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx51;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx52;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx53;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx54;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx56;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx57;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx58;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx60;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx61;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx62;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx63;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx65;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx66;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx67;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx69;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx72;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx73;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx76;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx78;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx80;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx82;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx83;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx84;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx87;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx91;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx92;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx95;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx102;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx103;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx105;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx109;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx110;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx114;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx117;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx118;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx120;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx122;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx123;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx127;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx128;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx131;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx134;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx135;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx136;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx138;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx140;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx146;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx147;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx148;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx149;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx152;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx153;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx156;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx157;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx158;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx159;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx160;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx162;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx163;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx168;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx170;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx171;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx172;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx173;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx175;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx177;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx178;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx181;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx182;
  wire multm_reduce_mulb0_add3b_maj3b_or3b_wx183;
  wire multm_reduce_mulb0_add3b_maj3b_wx2;
  wire multm_reduce_mulb0_add3b_maj3b_wx4;
  wire multm_reduce_mulb0_add3b_maj3b_wx8;
  wire multm_reduce_mulb0_add3b_maj3b_wx9;
  wire multm_reduce_mulb0_add3b_maj3b_wx12;
  wire multm_reduce_mulb0_add3b_maj3b_wx15;
  wire multm_reduce_mulb0_add3b_maj3b_wx16;
  wire multm_reduce_mulb0_add3b_maj3b_wx17;
  wire multm_reduce_mulb0_add3b_maj3b_wx18;
  wire multm_reduce_mulb0_add3b_maj3b_wx19;
  wire multm_reduce_mulb0_add3b_maj3b_wx20;
  wire multm_reduce_mulb0_add3b_maj3b_wx25;
  wire multm_reduce_mulb0_add3b_maj3b_wx26;
  wire multm_reduce_mulb0_add3b_maj3b_wx27;
  wire multm_reduce_mulb0_add3b_maj3b_wx29;
  wire multm_reduce_mulb0_add3b_maj3b_wx30;
  wire multm_reduce_mulb0_add3b_maj3b_wx33;
  wire multm_reduce_mulb0_add3b_maj3b_wx37;
  wire multm_reduce_mulb0_add3b_maj3b_wx40;
  wire multm_reduce_mulb0_add3b_maj3b_wx42;
  wire multm_reduce_mulb0_add3b_maj3b_wx44;
  wire multm_reduce_mulb0_add3b_maj3b_wx45;
  wire multm_reduce_mulb0_add3b_maj3b_wx46;
  wire multm_reduce_mulb0_add3b_maj3b_wx48;
  wire multm_reduce_mulb0_add3b_maj3b_wx50;
  wire multm_reduce_mulb0_add3b_maj3b_wx51;
  wire multm_reduce_mulb0_add3b_maj3b_wx52;
  wire multm_reduce_mulb0_add3b_maj3b_wx53;
  wire multm_reduce_mulb0_add3b_maj3b_wx54;
  wire multm_reduce_mulb0_add3b_maj3b_wx56;
  wire multm_reduce_mulb0_add3b_maj3b_wx57;
  wire multm_reduce_mulb0_add3b_maj3b_wx58;
  wire multm_reduce_mulb0_add3b_maj3b_wx60;
  wire multm_reduce_mulb0_add3b_maj3b_wx61;
  wire multm_reduce_mulb0_add3b_maj3b_wx62;
  wire multm_reduce_mulb0_add3b_maj3b_wx63;
  wire multm_reduce_mulb0_add3b_maj3b_wx65;
  wire multm_reduce_mulb0_add3b_maj3b_wx66;
  wire multm_reduce_mulb0_add3b_maj3b_wx67;
  wire multm_reduce_mulb0_add3b_maj3b_wx69;
  wire multm_reduce_mulb0_add3b_maj3b_wx72;
  wire multm_reduce_mulb0_add3b_maj3b_wx73;
  wire multm_reduce_mulb0_add3b_maj3b_wx76;
  wire multm_reduce_mulb0_add3b_maj3b_wx78;
  wire multm_reduce_mulb0_add3b_maj3b_wx80;
  wire multm_reduce_mulb0_add3b_maj3b_wx82;
  wire multm_reduce_mulb0_add3b_maj3b_wx83;
  wire multm_reduce_mulb0_add3b_maj3b_wx84;
  wire multm_reduce_mulb0_add3b_maj3b_wx87;
  wire multm_reduce_mulb0_add3b_maj3b_wx91;
  wire multm_reduce_mulb0_add3b_maj3b_wx92;
  wire multm_reduce_mulb0_add3b_maj3b_wx95;
  wire multm_reduce_mulb0_add3b_maj3b_wx102;
  wire multm_reduce_mulb0_add3b_maj3b_wx103;
  wire multm_reduce_mulb0_add3b_maj3b_wx105;
  wire multm_reduce_mulb0_add3b_maj3b_wx109;
  wire multm_reduce_mulb0_add3b_maj3b_wx110;
  wire multm_reduce_mulb0_add3b_maj3b_wx114;
  wire multm_reduce_mulb0_add3b_maj3b_wx117;
  wire multm_reduce_mulb0_add3b_maj3b_wx118;
  wire multm_reduce_mulb0_add3b_maj3b_wx120;
  wire multm_reduce_mulb0_add3b_maj3b_wx122;
  wire multm_reduce_mulb0_add3b_maj3b_wx123;
  wire multm_reduce_mulb0_add3b_maj3b_wx127;
  wire multm_reduce_mulb0_add3b_maj3b_wx128;
  wire multm_reduce_mulb0_add3b_maj3b_wx131;
  wire multm_reduce_mulb0_add3b_maj3b_wx134;
  wire multm_reduce_mulb0_add3b_maj3b_wx135;
  wire multm_reduce_mulb0_add3b_maj3b_wx136;
  wire multm_reduce_mulb0_add3b_maj3b_wx138;
  wire multm_reduce_mulb0_add3b_maj3b_wx140;
  wire multm_reduce_mulb0_add3b_maj3b_wx146;
  wire multm_reduce_mulb0_add3b_maj3b_wx147;
  wire multm_reduce_mulb0_add3b_maj3b_wx148;
  wire multm_reduce_mulb0_add3b_maj3b_wx149;
  wire multm_reduce_mulb0_add3b_maj3b_wx152;
  wire multm_reduce_mulb0_add3b_maj3b_wx153;
  wire multm_reduce_mulb0_add3b_maj3b_wx156;
  wire multm_reduce_mulb0_add3b_maj3b_wx157;
  wire multm_reduce_mulb0_add3b_maj3b_wx158;
  wire multm_reduce_mulb0_add3b_maj3b_wx159;
  wire multm_reduce_mulb0_add3b_maj3b_wx160;
  wire multm_reduce_mulb0_add3b_maj3b_wx162;
  wire multm_reduce_mulb0_add3b_maj3b_wx163;
  wire multm_reduce_mulb0_add3b_maj3b_wx168;
  wire multm_reduce_mulb0_add3b_maj3b_wx170;
  wire multm_reduce_mulb0_add3b_maj3b_wx171;
  wire multm_reduce_mulb0_add3b_maj3b_wx172;
  wire multm_reduce_mulb0_add3b_maj3b_wx173;
  wire multm_reduce_mulb0_add3b_maj3b_wx175;
  wire multm_reduce_mulb0_add3b_maj3b_wx177;
  wire multm_reduce_mulb0_add3b_maj3b_wx178;
  wire multm_reduce_mulb0_add3b_maj3b_wx181;
  wire multm_reduce_mulb0_add3b_maj3b_wx182;
  wire multm_reduce_mulb0_add3b_maj3b_wx183;
  wire multm_reduce_mulb0_add3b_maj3b_wy2;
  wire multm_reduce_mulb0_add3b_maj3b_wy4;
  wire multm_reduce_mulb0_add3b_maj3b_wy8;
  wire multm_reduce_mulb0_add3b_maj3b_wy9;
  wire multm_reduce_mulb0_add3b_maj3b_wy12;
  wire multm_reduce_mulb0_add3b_maj3b_wy15;
  wire multm_reduce_mulb0_add3b_maj3b_wy16;
  wire multm_reduce_mulb0_add3b_maj3b_wy17;
  wire multm_reduce_mulb0_add3b_maj3b_wy18;
  wire multm_reduce_mulb0_add3b_maj3b_wy19;
  wire multm_reduce_mulb0_add3b_maj3b_wy20;
  wire multm_reduce_mulb0_add3b_maj3b_wy25;
  wire multm_reduce_mulb0_add3b_maj3b_wy26;
  wire multm_reduce_mulb0_add3b_maj3b_wy27;
  wire multm_reduce_mulb0_add3b_maj3b_wy29;
  wire multm_reduce_mulb0_add3b_maj3b_wy30;
  wire multm_reduce_mulb0_add3b_maj3b_wy33;
  wire multm_reduce_mulb0_add3b_maj3b_wy37;
  wire multm_reduce_mulb0_add3b_maj3b_wy40;
  wire multm_reduce_mulb0_add3b_maj3b_wy42;
  wire multm_reduce_mulb0_add3b_maj3b_wy44;
  wire multm_reduce_mulb0_add3b_maj3b_wy45;
  wire multm_reduce_mulb0_add3b_maj3b_wy46;
  wire multm_reduce_mulb0_add3b_maj3b_wy48;
  wire multm_reduce_mulb0_add3b_maj3b_wy50;
  wire multm_reduce_mulb0_add3b_maj3b_wy51;
  wire multm_reduce_mulb0_add3b_maj3b_wy52;
  wire multm_reduce_mulb0_add3b_maj3b_wy53;
  wire multm_reduce_mulb0_add3b_maj3b_wy54;
  wire multm_reduce_mulb0_add3b_maj3b_wy56;
  wire multm_reduce_mulb0_add3b_maj3b_wy57;
  wire multm_reduce_mulb0_add3b_maj3b_wy58;
  wire multm_reduce_mulb0_add3b_maj3b_wy60;
  wire multm_reduce_mulb0_add3b_maj3b_wy61;
  wire multm_reduce_mulb0_add3b_maj3b_wy62;
  wire multm_reduce_mulb0_add3b_maj3b_wy63;
  wire multm_reduce_mulb0_add3b_maj3b_wy65;
  wire multm_reduce_mulb0_add3b_maj3b_wy66;
  wire multm_reduce_mulb0_add3b_maj3b_wy67;
  wire multm_reduce_mulb0_add3b_maj3b_wy69;
  wire multm_reduce_mulb0_add3b_maj3b_wy72;
  wire multm_reduce_mulb0_add3b_maj3b_wy73;
  wire multm_reduce_mulb0_add3b_maj3b_wy76;
  wire multm_reduce_mulb0_add3b_maj3b_wy78;
  wire multm_reduce_mulb0_add3b_maj3b_wy80;
  wire multm_reduce_mulb0_add3b_maj3b_wy82;
  wire multm_reduce_mulb0_add3b_maj3b_wy83;
  wire multm_reduce_mulb0_add3b_maj3b_wy84;
  wire multm_reduce_mulb0_add3b_maj3b_wy87;
  wire multm_reduce_mulb0_add3b_maj3b_wy91;
  wire multm_reduce_mulb0_add3b_maj3b_wy92;
  wire multm_reduce_mulb0_add3b_maj3b_wy95;
  wire multm_reduce_mulb0_add3b_maj3b_wy102;
  wire multm_reduce_mulb0_add3b_maj3b_wy103;
  wire multm_reduce_mulb0_add3b_maj3b_wy105;
  wire multm_reduce_mulb0_add3b_maj3b_wy109;
  wire multm_reduce_mulb0_add3b_maj3b_wy110;
  wire multm_reduce_mulb0_add3b_maj3b_wy114;
  wire multm_reduce_mulb0_add3b_maj3b_wy117;
  wire multm_reduce_mulb0_add3b_maj3b_wy118;
  wire multm_reduce_mulb0_add3b_maj3b_wy120;
  wire multm_reduce_mulb0_add3b_maj3b_wy122;
  wire multm_reduce_mulb0_add3b_maj3b_wy123;
  wire multm_reduce_mulb0_add3b_maj3b_wy127;
  wire multm_reduce_mulb0_add3b_maj3b_wy128;
  wire multm_reduce_mulb0_add3b_maj3b_wy131;
  wire multm_reduce_mulb0_add3b_maj3b_wy134;
  wire multm_reduce_mulb0_add3b_maj3b_wy135;
  wire multm_reduce_mulb0_add3b_maj3b_wy136;
  wire multm_reduce_mulb0_add3b_maj3b_wy138;
  wire multm_reduce_mulb0_add3b_maj3b_wy140;
  wire multm_reduce_mulb0_add3b_maj3b_wy146;
  wire multm_reduce_mulb0_add3b_maj3b_wy147;
  wire multm_reduce_mulb0_add3b_maj3b_wy148;
  wire multm_reduce_mulb0_add3b_maj3b_wy149;
  wire multm_reduce_mulb0_add3b_maj3b_wy152;
  wire multm_reduce_mulb0_add3b_maj3b_wy153;
  wire multm_reduce_mulb0_add3b_maj3b_wy156;
  wire multm_reduce_mulb0_add3b_maj3b_wy157;
  wire multm_reduce_mulb0_add3b_maj3b_wy158;
  wire multm_reduce_mulb0_add3b_maj3b_wy159;
  wire multm_reduce_mulb0_add3b_maj3b_wy160;
  wire multm_reduce_mulb0_add3b_maj3b_wy162;
  wire multm_reduce_mulb0_add3b_maj3b_wy163;
  wire multm_reduce_mulb0_add3b_maj3b_wy168;
  wire multm_reduce_mulb0_add3b_maj3b_wy170;
  wire multm_reduce_mulb0_add3b_maj3b_wy171;
  wire multm_reduce_mulb0_add3b_maj3b_wy172;
  wire multm_reduce_mulb0_add3b_maj3b_wy173;
  wire multm_reduce_mulb0_add3b_maj3b_wy175;
  wire multm_reduce_mulb0_add3b_maj3b_wy177;
  wire multm_reduce_mulb0_add3b_maj3b_wy178;
  wire multm_reduce_mulb0_add3b_maj3b_wy181;
  wire multm_reduce_mulb0_add3b_maj3b_wy182;
  wire multm_reduce_mulb0_add3b_maj3b_wy183;
  wire multm_reduce_mulb0_add3b_maj3b_xy2;
  wire multm_reduce_mulb0_add3b_maj3b_xy4;
  wire multm_reduce_mulb0_add3b_maj3b_xy8;
  wire multm_reduce_mulb0_add3b_maj3b_xy9;
  wire multm_reduce_mulb0_add3b_maj3b_xy12;
  wire multm_reduce_mulb0_add3b_maj3b_xy15;
  wire multm_reduce_mulb0_add3b_maj3b_xy16;
  wire multm_reduce_mulb0_add3b_maj3b_xy17;
  wire multm_reduce_mulb0_add3b_maj3b_xy18;
  wire multm_reduce_mulb0_add3b_maj3b_xy19;
  wire multm_reduce_mulb0_add3b_maj3b_xy20;
  wire multm_reduce_mulb0_add3b_maj3b_xy25;
  wire multm_reduce_mulb0_add3b_maj3b_xy26;
  wire multm_reduce_mulb0_add3b_maj3b_xy27;
  wire multm_reduce_mulb0_add3b_maj3b_xy29;
  wire multm_reduce_mulb0_add3b_maj3b_xy30;
  wire multm_reduce_mulb0_add3b_maj3b_xy33;
  wire multm_reduce_mulb0_add3b_maj3b_xy37;
  wire multm_reduce_mulb0_add3b_maj3b_xy40;
  wire multm_reduce_mulb0_add3b_maj3b_xy42;
  wire multm_reduce_mulb0_add3b_maj3b_xy44;
  wire multm_reduce_mulb0_add3b_maj3b_xy45;
  wire multm_reduce_mulb0_add3b_maj3b_xy46;
  wire multm_reduce_mulb0_add3b_maj3b_xy48;
  wire multm_reduce_mulb0_add3b_maj3b_xy50;
  wire multm_reduce_mulb0_add3b_maj3b_xy51;
  wire multm_reduce_mulb0_add3b_maj3b_xy52;
  wire multm_reduce_mulb0_add3b_maj3b_xy53;
  wire multm_reduce_mulb0_add3b_maj3b_xy54;
  wire multm_reduce_mulb0_add3b_maj3b_xy56;
  wire multm_reduce_mulb0_add3b_maj3b_xy57;
  wire multm_reduce_mulb0_add3b_maj3b_xy58;
  wire multm_reduce_mulb0_add3b_maj3b_xy60;
  wire multm_reduce_mulb0_add3b_maj3b_xy61;
  wire multm_reduce_mulb0_add3b_maj3b_xy62;
  wire multm_reduce_mulb0_add3b_maj3b_xy63;
  wire multm_reduce_mulb0_add3b_maj3b_xy65;
  wire multm_reduce_mulb0_add3b_maj3b_xy66;
  wire multm_reduce_mulb0_add3b_maj3b_xy67;
  wire multm_reduce_mulb0_add3b_maj3b_xy69;
  wire multm_reduce_mulb0_add3b_maj3b_xy72;
  wire multm_reduce_mulb0_add3b_maj3b_xy73;
  wire multm_reduce_mulb0_add3b_maj3b_xy76;
  wire multm_reduce_mulb0_add3b_maj3b_xy78;
  wire multm_reduce_mulb0_add3b_maj3b_xy80;
  wire multm_reduce_mulb0_add3b_maj3b_xy82;
  wire multm_reduce_mulb0_add3b_maj3b_xy83;
  wire multm_reduce_mulb0_add3b_maj3b_xy84;
  wire multm_reduce_mulb0_add3b_maj3b_xy87;
  wire multm_reduce_mulb0_add3b_maj3b_xy91;
  wire multm_reduce_mulb0_add3b_maj3b_xy92;
  wire multm_reduce_mulb0_add3b_maj3b_xy95;
  wire multm_reduce_mulb0_add3b_maj3b_xy102;
  wire multm_reduce_mulb0_add3b_maj3b_xy103;
  wire multm_reduce_mulb0_add3b_maj3b_xy105;
  wire multm_reduce_mulb0_add3b_maj3b_xy109;
  wire multm_reduce_mulb0_add3b_maj3b_xy110;
  wire multm_reduce_mulb0_add3b_maj3b_xy114;
  wire multm_reduce_mulb0_add3b_maj3b_xy117;
  wire multm_reduce_mulb0_add3b_maj3b_xy118;
  wire multm_reduce_mulb0_add3b_maj3b_xy120;
  wire multm_reduce_mulb0_add3b_maj3b_xy122;
  wire multm_reduce_mulb0_add3b_maj3b_xy123;
  wire multm_reduce_mulb0_add3b_maj3b_xy127;
  wire multm_reduce_mulb0_add3b_maj3b_xy128;
  wire multm_reduce_mulb0_add3b_maj3b_xy131;
  wire multm_reduce_mulb0_add3b_maj3b_xy134;
  wire multm_reduce_mulb0_add3b_maj3b_xy135;
  wire multm_reduce_mulb0_add3b_maj3b_xy136;
  wire multm_reduce_mulb0_add3b_maj3b_xy138;
  wire multm_reduce_mulb0_add3b_maj3b_xy140;
  wire multm_reduce_mulb0_add3b_maj3b_xy146;
  wire multm_reduce_mulb0_add3b_maj3b_xy147;
  wire multm_reduce_mulb0_add3b_maj3b_xy148;
  wire multm_reduce_mulb0_add3b_maj3b_xy149;
  wire multm_reduce_mulb0_add3b_maj3b_xy152;
  wire multm_reduce_mulb0_add3b_maj3b_xy153;
  wire multm_reduce_mulb0_add3b_maj3b_xy156;
  wire multm_reduce_mulb0_add3b_maj3b_xy157;
  wire multm_reduce_mulb0_add3b_maj3b_xy158;
  wire multm_reduce_mulb0_add3b_maj3b_xy159;
  wire multm_reduce_mulb0_add3b_maj3b_xy160;
  wire multm_reduce_mulb0_add3b_maj3b_xy162;
  wire multm_reduce_mulb0_add3b_maj3b_xy163;
  wire multm_reduce_mulb0_add3b_maj3b_xy168;
  wire multm_reduce_mulb0_add3b_maj3b_xy170;
  wire multm_reduce_mulb0_add3b_maj3b_xy171;
  wire multm_reduce_mulb0_add3b_maj3b_xy172;
  wire multm_reduce_mulb0_add3b_maj3b_xy173;
  wire multm_reduce_mulb0_add3b_maj3b_xy175;
  wire multm_reduce_mulb0_add3b_maj3b_xy177;
  wire multm_reduce_mulb0_add3b_maj3b_xy178;
  wire multm_reduce_mulb0_add3b_maj3b_xy181;
  wire multm_reduce_mulb0_add3b_maj3b_xy182;
  wire multm_reduce_mulb0_add3b_maj3b_xy183;
  wire multm_reduce_mulb0_add3b_xor3b_wx2;
  wire multm_reduce_mulb0_add3b_xor3b_wx4;
  wire multm_reduce_mulb0_add3b_xor3b_wx8;
  wire multm_reduce_mulb0_add3b_xor3b_wx9;
  wire multm_reduce_mulb0_add3b_xor3b_wx12;
  wire multm_reduce_mulb0_add3b_xor3b_wx15;
  wire multm_reduce_mulb0_add3b_xor3b_wx16;
  wire multm_reduce_mulb0_add3b_xor3b_wx17;
  wire multm_reduce_mulb0_add3b_xor3b_wx18;
  wire multm_reduce_mulb0_add3b_xor3b_wx19;
  wire multm_reduce_mulb0_add3b_xor3b_wx20;
  wire multm_reduce_mulb0_add3b_xor3b_wx25;
  wire multm_reduce_mulb0_add3b_xor3b_wx26;
  wire multm_reduce_mulb0_add3b_xor3b_wx27;
  wire multm_reduce_mulb0_add3b_xor3b_wx29;
  wire multm_reduce_mulb0_add3b_xor3b_wx30;
  wire multm_reduce_mulb0_add3b_xor3b_wx33;
  wire multm_reduce_mulb0_add3b_xor3b_wx37;
  wire multm_reduce_mulb0_add3b_xor3b_wx40;
  wire multm_reduce_mulb0_add3b_xor3b_wx42;
  wire multm_reduce_mulb0_add3b_xor3b_wx44;
  wire multm_reduce_mulb0_add3b_xor3b_wx45;
  wire multm_reduce_mulb0_add3b_xor3b_wx46;
  wire multm_reduce_mulb0_add3b_xor3b_wx48;
  wire multm_reduce_mulb0_add3b_xor3b_wx50;
  wire multm_reduce_mulb0_add3b_xor3b_wx51;
  wire multm_reduce_mulb0_add3b_xor3b_wx52;
  wire multm_reduce_mulb0_add3b_xor3b_wx53;
  wire multm_reduce_mulb0_add3b_xor3b_wx54;
  wire multm_reduce_mulb0_add3b_xor3b_wx56;
  wire multm_reduce_mulb0_add3b_xor3b_wx57;
  wire multm_reduce_mulb0_add3b_xor3b_wx58;
  wire multm_reduce_mulb0_add3b_xor3b_wx60;
  wire multm_reduce_mulb0_add3b_xor3b_wx61;
  wire multm_reduce_mulb0_add3b_xor3b_wx62;
  wire multm_reduce_mulb0_add3b_xor3b_wx63;
  wire multm_reduce_mulb0_add3b_xor3b_wx65;
  wire multm_reduce_mulb0_add3b_xor3b_wx66;
  wire multm_reduce_mulb0_add3b_xor3b_wx67;
  wire multm_reduce_mulb0_add3b_xor3b_wx69;
  wire multm_reduce_mulb0_add3b_xor3b_wx72;
  wire multm_reduce_mulb0_add3b_xor3b_wx73;
  wire multm_reduce_mulb0_add3b_xor3b_wx76;
  wire multm_reduce_mulb0_add3b_xor3b_wx78;
  wire multm_reduce_mulb0_add3b_xor3b_wx80;
  wire multm_reduce_mulb0_add3b_xor3b_wx82;
  wire multm_reduce_mulb0_add3b_xor3b_wx83;
  wire multm_reduce_mulb0_add3b_xor3b_wx84;
  wire multm_reduce_mulb0_add3b_xor3b_wx87;
  wire multm_reduce_mulb0_add3b_xor3b_wx91;
  wire multm_reduce_mulb0_add3b_xor3b_wx92;
  wire multm_reduce_mulb0_add3b_xor3b_wx95;
  wire multm_reduce_mulb0_add3b_xor3b_wx102;
  wire multm_reduce_mulb0_add3b_xor3b_wx103;
  wire multm_reduce_mulb0_add3b_xor3b_wx105;
  wire multm_reduce_mulb0_add3b_xor3b_wx109;
  wire multm_reduce_mulb0_add3b_xor3b_wx110;
  wire multm_reduce_mulb0_add3b_xor3b_wx114;
  wire multm_reduce_mulb0_add3b_xor3b_wx117;
  wire multm_reduce_mulb0_add3b_xor3b_wx118;
  wire multm_reduce_mulb0_add3b_xor3b_wx120;
  wire multm_reduce_mulb0_add3b_xor3b_wx122;
  wire multm_reduce_mulb0_add3b_xor3b_wx123;
  wire multm_reduce_mulb0_add3b_xor3b_wx127;
  wire multm_reduce_mulb0_add3b_xor3b_wx128;
  wire multm_reduce_mulb0_add3b_xor3b_wx131;
  wire multm_reduce_mulb0_add3b_xor3b_wx134;
  wire multm_reduce_mulb0_add3b_xor3b_wx135;
  wire multm_reduce_mulb0_add3b_xor3b_wx136;
  wire multm_reduce_mulb0_add3b_xor3b_wx138;
  wire multm_reduce_mulb0_add3b_xor3b_wx140;
  wire multm_reduce_mulb0_add3b_xor3b_wx146;
  wire multm_reduce_mulb0_add3b_xor3b_wx147;
  wire multm_reduce_mulb0_add3b_xor3b_wx148;
  wire multm_reduce_mulb0_add3b_xor3b_wx149;
  wire multm_reduce_mulb0_add3b_xor3b_wx152;
  wire multm_reduce_mulb0_add3b_xor3b_wx153;
  wire multm_reduce_mulb0_add3b_xor3b_wx156;
  wire multm_reduce_mulb0_add3b_xor3b_wx157;
  wire multm_reduce_mulb0_add3b_xor3b_wx158;
  wire multm_reduce_mulb0_add3b_xor3b_wx159;
  wire multm_reduce_mulb0_add3b_xor3b_wx160;
  wire multm_reduce_mulb0_add3b_xor3b_wx162;
  wire multm_reduce_mulb0_add3b_xor3b_wx163;
  wire multm_reduce_mulb0_add3b_xor3b_wx168;
  wire multm_reduce_mulb0_add3b_xor3b_wx170;
  wire multm_reduce_mulb0_add3b_xor3b_wx171;
  wire multm_reduce_mulb0_add3b_xor3b_wx172;
  wire multm_reduce_mulb0_add3b_xor3b_wx173;
  wire multm_reduce_mulb0_add3b_xor3b_wx175;
  wire multm_reduce_mulb0_add3b_xor3b_wx177;
  wire multm_reduce_mulb0_add3b_xor3b_wx178;
  wire multm_reduce_mulb0_add3b_xor3b_wx181;
  wire multm_reduce_mulb0_add3b_xor3b_wx182;
  wire multm_reduce_mulb0_add3b_xor3b_wx183;
  wire multm_reduce_mulb0_cq0;
  wire multm_reduce_mulb0_cq1;
  wire multm_reduce_mulb0_cq2;
  wire multm_reduce_mulb0_cq3;
  wire multm_reduce_mulb0_cq4;
  wire multm_reduce_mulb0_cq5;
  wire multm_reduce_mulb0_cq6;
  wire multm_reduce_mulb0_cq7;
  wire multm_reduce_mulb0_cq8;
  wire multm_reduce_mulb0_cq9;
  wire multm_reduce_mulb0_cq10;
  wire multm_reduce_mulb0_cq11;
  wire multm_reduce_mulb0_cq12;
  wire multm_reduce_mulb0_cq13;
  wire multm_reduce_mulb0_cq14;
  wire multm_reduce_mulb0_cq15;
  wire multm_reduce_mulb0_cq16;
  wire multm_reduce_mulb0_cq17;
  wire multm_reduce_mulb0_cq18;
  wire multm_reduce_mulb0_cq19;
  wire multm_reduce_mulb0_cq20;
  wire multm_reduce_mulb0_cq21;
  wire multm_reduce_mulb0_cq22;
  wire multm_reduce_mulb0_cq23;
  wire multm_reduce_mulb0_cq24;
  wire multm_reduce_mulb0_cq25;
  wire multm_reduce_mulb0_cq26;
  wire multm_reduce_mulb0_cq27;
  wire multm_reduce_mulb0_cq28;
  wire multm_reduce_mulb0_cq29;
  wire multm_reduce_mulb0_cq30;
  wire multm_reduce_mulb0_cq31;
  wire multm_reduce_mulb0_cq32;
  wire multm_reduce_mulb0_cq33;
  wire multm_reduce_mulb0_cq34;
  wire multm_reduce_mulb0_cq35;
  wire multm_reduce_mulb0_cq36;
  wire multm_reduce_mulb0_cq37;
  wire multm_reduce_mulb0_cq38;
  wire multm_reduce_mulb0_cq39;
  wire multm_reduce_mulb0_cq40;
  wire multm_reduce_mulb0_cq41;
  wire multm_reduce_mulb0_cq42;
  wire multm_reduce_mulb0_cq43;
  wire multm_reduce_mulb0_cq44;
  wire multm_reduce_mulb0_cq45;
  wire multm_reduce_mulb0_cq46;
  wire multm_reduce_mulb0_cq47;
  wire multm_reduce_mulb0_cq48;
  wire multm_reduce_mulb0_cq49;
  wire multm_reduce_mulb0_cq50;
  wire multm_reduce_mulb0_cq51;
  wire multm_reduce_mulb0_cq52;
  wire multm_reduce_mulb0_cq53;
  wire multm_reduce_mulb0_cq54;
  wire multm_reduce_mulb0_cq55;
  wire multm_reduce_mulb0_cq56;
  wire multm_reduce_mulb0_cq57;
  wire multm_reduce_mulb0_cq58;
  wire multm_reduce_mulb0_cq59;
  wire multm_reduce_mulb0_cq60;
  wire multm_reduce_mulb0_cq61;
  wire multm_reduce_mulb0_cq62;
  wire multm_reduce_mulb0_cq63;
  wire multm_reduce_mulb0_cq64;
  wire multm_reduce_mulb0_cq65;
  wire multm_reduce_mulb0_cq66;
  wire multm_reduce_mulb0_cq67;
  wire multm_reduce_mulb0_cq68;
  wire multm_reduce_mulb0_cq69;
  wire multm_reduce_mulb0_cq70;
  wire multm_reduce_mulb0_cq71;
  wire multm_reduce_mulb0_cq72;
  wire multm_reduce_mulb0_cq73;
  wire multm_reduce_mulb0_cq74;
  wire multm_reduce_mulb0_cq75;
  wire multm_reduce_mulb0_cq76;
  wire multm_reduce_mulb0_cq77;
  wire multm_reduce_mulb0_cq78;
  wire multm_reduce_mulb0_cq79;
  wire multm_reduce_mulb0_cq80;
  wire multm_reduce_mulb0_cq81;
  wire multm_reduce_mulb0_cq82;
  wire multm_reduce_mulb0_cq83;
  wire multm_reduce_mulb0_cq84;
  wire multm_reduce_mulb0_cq85;
  wire multm_reduce_mulb0_cq86;
  wire multm_reduce_mulb0_cq87;
  wire multm_reduce_mulb0_cq88;
  wire multm_reduce_mulb0_cq89;
  wire multm_reduce_mulb0_cq90;
  wire multm_reduce_mulb0_cq91;
  wire multm_reduce_mulb0_cq92;
  wire multm_reduce_mulb0_cq93;
  wire multm_reduce_mulb0_cq94;
  wire multm_reduce_mulb0_cq95;
  wire multm_reduce_mulb0_cq96;
  wire multm_reduce_mulb0_cq97;
  wire multm_reduce_mulb0_cq98;
  wire multm_reduce_mulb0_cq99;
  wire multm_reduce_mulb0_cq100;
  wire multm_reduce_mulb0_cq101;
  wire multm_reduce_mulb0_cq102;
  wire multm_reduce_mulb0_cq103;
  wire multm_reduce_mulb0_cq104;
  wire multm_reduce_mulb0_cq105;
  wire multm_reduce_mulb0_cq106;
  wire multm_reduce_mulb0_cq107;
  wire multm_reduce_mulb0_cq108;
  wire multm_reduce_mulb0_cq109;
  wire multm_reduce_mulb0_cq110;
  wire multm_reduce_mulb0_cq111;
  wire multm_reduce_mulb0_cq112;
  wire multm_reduce_mulb0_cq113;
  wire multm_reduce_mulb0_cq114;
  wire multm_reduce_mulb0_cq115;
  wire multm_reduce_mulb0_cq116;
  wire multm_reduce_mulb0_cq117;
  wire multm_reduce_mulb0_cq118;
  wire multm_reduce_mulb0_cq119;
  wire multm_reduce_mulb0_cq120;
  wire multm_reduce_mulb0_cq121;
  wire multm_reduce_mulb0_cq122;
  wire multm_reduce_mulb0_cq123;
  wire multm_reduce_mulb0_cq124;
  wire multm_reduce_mulb0_cq125;
  wire multm_reduce_mulb0_cq126;
  wire multm_reduce_mulb0_cq127;
  wire multm_reduce_mulb0_cq128;
  wire multm_reduce_mulb0_cq129;
  wire multm_reduce_mulb0_cq130;
  wire multm_reduce_mulb0_cq131;
  wire multm_reduce_mulb0_cq132;
  wire multm_reduce_mulb0_cq133;
  wire multm_reduce_mulb0_cq134;
  wire multm_reduce_mulb0_cq135;
  wire multm_reduce_mulb0_cq136;
  wire multm_reduce_mulb0_cq137;
  wire multm_reduce_mulb0_cq138;
  wire multm_reduce_mulb0_cq139;
  wire multm_reduce_mulb0_cq140;
  wire multm_reduce_mulb0_cq141;
  wire multm_reduce_mulb0_cq142;
  wire multm_reduce_mulb0_cq143;
  wire multm_reduce_mulb0_cq144;
  wire multm_reduce_mulb0_cq145;
  wire multm_reduce_mulb0_cq146;
  wire multm_reduce_mulb0_cq147;
  wire multm_reduce_mulb0_cq148;
  wire multm_reduce_mulb0_cq149;
  wire multm_reduce_mulb0_cq150;
  wire multm_reduce_mulb0_cq151;
  wire multm_reduce_mulb0_cq152;
  wire multm_reduce_mulb0_cq153;
  wire multm_reduce_mulb0_cq154;
  wire multm_reduce_mulb0_cq155;
  wire multm_reduce_mulb0_cq156;
  wire multm_reduce_mulb0_cq157;
  wire multm_reduce_mulb0_cq158;
  wire multm_reduce_mulb0_cq159;
  wire multm_reduce_mulb0_cq160;
  wire multm_reduce_mulb0_cq161;
  wire multm_reduce_mulb0_cq162;
  wire multm_reduce_mulb0_cq163;
  wire multm_reduce_mulb0_cq164;
  wire multm_reduce_mulb0_cq165;
  wire multm_reduce_mulb0_cq166;
  wire multm_reduce_mulb0_cq167;
  wire multm_reduce_mulb0_cq168;
  wire multm_reduce_mulb0_cq169;
  wire multm_reduce_mulb0_cq170;
  wire multm_reduce_mulb0_cq171;
  wire multm_reduce_mulb0_cq172;
  wire multm_reduce_mulb0_cq173;
  wire multm_reduce_mulb0_cq174;
  wire multm_reduce_mulb0_cq175;
  wire multm_reduce_mulb0_cq176;
  wire multm_reduce_mulb0_cq177;
  wire multm_reduce_mulb0_cq178;
  wire multm_reduce_mulb0_cq179;
  wire multm_reduce_mulb0_cq180;
  wire multm_reduce_mulb0_cq181;
  wire multm_reduce_mulb0_cq182;
  wire multm_reduce_mulb0_cq183;
  wire multm_reduce_mulb0_cq184;
  wire multm_reduce_mulb0_pc0;
  wire multm_reduce_mulb0_pc1;
  wire multm_reduce_mulb0_pc2;
  wire multm_reduce_mulb0_pc3;
  wire multm_reduce_mulb0_pc4;
  wire multm_reduce_mulb0_pc5;
  wire multm_reduce_mulb0_pc6;
  wire multm_reduce_mulb0_pc7;
  wire multm_reduce_mulb0_pc8;
  wire multm_reduce_mulb0_pc9;
  wire multm_reduce_mulb0_pc10;
  wire multm_reduce_mulb0_pc11;
  wire multm_reduce_mulb0_pc12;
  wire multm_reduce_mulb0_pc13;
  wire multm_reduce_mulb0_pc14;
  wire multm_reduce_mulb0_pc15;
  wire multm_reduce_mulb0_pc16;
  wire multm_reduce_mulb0_pc17;
  wire multm_reduce_mulb0_pc18;
  wire multm_reduce_mulb0_pc19;
  wire multm_reduce_mulb0_pc20;
  wire multm_reduce_mulb0_pc21;
  wire multm_reduce_mulb0_pc22;
  wire multm_reduce_mulb0_pc23;
  wire multm_reduce_mulb0_pc24;
  wire multm_reduce_mulb0_pc25;
  wire multm_reduce_mulb0_pc26;
  wire multm_reduce_mulb0_pc27;
  wire multm_reduce_mulb0_pc28;
  wire multm_reduce_mulb0_pc29;
  wire multm_reduce_mulb0_pc30;
  wire multm_reduce_mulb0_pc31;
  wire multm_reduce_mulb0_pc32;
  wire multm_reduce_mulb0_pc33;
  wire multm_reduce_mulb0_pc34;
  wire multm_reduce_mulb0_pc35;
  wire multm_reduce_mulb0_pc36;
  wire multm_reduce_mulb0_pc37;
  wire multm_reduce_mulb0_pc38;
  wire multm_reduce_mulb0_pc39;
  wire multm_reduce_mulb0_pc40;
  wire multm_reduce_mulb0_pc41;
  wire multm_reduce_mulb0_pc42;
  wire multm_reduce_mulb0_pc43;
  wire multm_reduce_mulb0_pc44;
  wire multm_reduce_mulb0_pc45;
  wire multm_reduce_mulb0_pc46;
  wire multm_reduce_mulb0_pc47;
  wire multm_reduce_mulb0_pc48;
  wire multm_reduce_mulb0_pc49;
  wire multm_reduce_mulb0_pc50;
  wire multm_reduce_mulb0_pc51;
  wire multm_reduce_mulb0_pc52;
  wire multm_reduce_mulb0_pc53;
  wire multm_reduce_mulb0_pc54;
  wire multm_reduce_mulb0_pc55;
  wire multm_reduce_mulb0_pc56;
  wire multm_reduce_mulb0_pc57;
  wire multm_reduce_mulb0_pc58;
  wire multm_reduce_mulb0_pc59;
  wire multm_reduce_mulb0_pc60;
  wire multm_reduce_mulb0_pc61;
  wire multm_reduce_mulb0_pc62;
  wire multm_reduce_mulb0_pc63;
  wire multm_reduce_mulb0_pc64;
  wire multm_reduce_mulb0_pc65;
  wire multm_reduce_mulb0_pc66;
  wire multm_reduce_mulb0_pc67;
  wire multm_reduce_mulb0_pc68;
  wire multm_reduce_mulb0_pc69;
  wire multm_reduce_mulb0_pc70;
  wire multm_reduce_mulb0_pc71;
  wire multm_reduce_mulb0_pc72;
  wire multm_reduce_mulb0_pc73;
  wire multm_reduce_mulb0_pc74;
  wire multm_reduce_mulb0_pc75;
  wire multm_reduce_mulb0_pc76;
  wire multm_reduce_mulb0_pc77;
  wire multm_reduce_mulb0_pc78;
  wire multm_reduce_mulb0_pc79;
  wire multm_reduce_mulb0_pc80;
  wire multm_reduce_mulb0_pc81;
  wire multm_reduce_mulb0_pc82;
  wire multm_reduce_mulb0_pc83;
  wire multm_reduce_mulb0_pc84;
  wire multm_reduce_mulb0_pc85;
  wire multm_reduce_mulb0_pc86;
  wire multm_reduce_mulb0_pc87;
  wire multm_reduce_mulb0_pc88;
  wire multm_reduce_mulb0_pc89;
  wire multm_reduce_mulb0_pc90;
  wire multm_reduce_mulb0_pc91;
  wire multm_reduce_mulb0_pc92;
  wire multm_reduce_mulb0_pc93;
  wire multm_reduce_mulb0_pc94;
  wire multm_reduce_mulb0_pc95;
  wire multm_reduce_mulb0_pc96;
  wire multm_reduce_mulb0_pc97;
  wire multm_reduce_mulb0_pc98;
  wire multm_reduce_mulb0_pc99;
  wire multm_reduce_mulb0_pc100;
  wire multm_reduce_mulb0_pc101;
  wire multm_reduce_mulb0_pc102;
  wire multm_reduce_mulb0_pc103;
  wire multm_reduce_mulb0_pc104;
  wire multm_reduce_mulb0_pc105;
  wire multm_reduce_mulb0_pc106;
  wire multm_reduce_mulb0_pc107;
  wire multm_reduce_mulb0_pc108;
  wire multm_reduce_mulb0_pc109;
  wire multm_reduce_mulb0_pc110;
  wire multm_reduce_mulb0_pc111;
  wire multm_reduce_mulb0_pc112;
  wire multm_reduce_mulb0_pc113;
  wire multm_reduce_mulb0_pc114;
  wire multm_reduce_mulb0_pc115;
  wire multm_reduce_mulb0_pc116;
  wire multm_reduce_mulb0_pc117;
  wire multm_reduce_mulb0_pc118;
  wire multm_reduce_mulb0_pc119;
  wire multm_reduce_mulb0_pc120;
  wire multm_reduce_mulb0_pc121;
  wire multm_reduce_mulb0_pc122;
  wire multm_reduce_mulb0_pc123;
  wire multm_reduce_mulb0_pc124;
  wire multm_reduce_mulb0_pc125;
  wire multm_reduce_mulb0_pc126;
  wire multm_reduce_mulb0_pc127;
  wire multm_reduce_mulb0_pc128;
  wire multm_reduce_mulb0_pc129;
  wire multm_reduce_mulb0_pc130;
  wire multm_reduce_mulb0_pc131;
  wire multm_reduce_mulb0_pc132;
  wire multm_reduce_mulb0_pc133;
  wire multm_reduce_mulb0_pc134;
  wire multm_reduce_mulb0_pc135;
  wire multm_reduce_mulb0_pc136;
  wire multm_reduce_mulb0_pc137;
  wire multm_reduce_mulb0_pc138;
  wire multm_reduce_mulb0_pc139;
  wire multm_reduce_mulb0_pc140;
  wire multm_reduce_mulb0_pc141;
  wire multm_reduce_mulb0_pc142;
  wire multm_reduce_mulb0_pc143;
  wire multm_reduce_mulb0_pc144;
  wire multm_reduce_mulb0_pc145;
  wire multm_reduce_mulb0_pc146;
  wire multm_reduce_mulb0_pc147;
  wire multm_reduce_mulb0_pc148;
  wire multm_reduce_mulb0_pc149;
  wire multm_reduce_mulb0_pc150;
  wire multm_reduce_mulb0_pc151;
  wire multm_reduce_mulb0_pc152;
  wire multm_reduce_mulb0_pc153;
  wire multm_reduce_mulb0_pc154;
  wire multm_reduce_mulb0_pc155;
  wire multm_reduce_mulb0_pc156;
  wire multm_reduce_mulb0_pc157;
  wire multm_reduce_mulb0_pc158;
  wire multm_reduce_mulb0_pc159;
  wire multm_reduce_mulb0_pc160;
  wire multm_reduce_mulb0_pc161;
  wire multm_reduce_mulb0_pc162;
  wire multm_reduce_mulb0_pc163;
  wire multm_reduce_mulb0_pc164;
  wire multm_reduce_mulb0_pc165;
  wire multm_reduce_mulb0_pc166;
  wire multm_reduce_mulb0_pc167;
  wire multm_reduce_mulb0_pc168;
  wire multm_reduce_mulb0_pc169;
  wire multm_reduce_mulb0_pc170;
  wire multm_reduce_mulb0_pc171;
  wire multm_reduce_mulb0_pc172;
  wire multm_reduce_mulb0_pc173;
  wire multm_reduce_mulb0_pc174;
  wire multm_reduce_mulb0_pc175;
  wire multm_reduce_mulb0_pc176;
  wire multm_reduce_mulb0_pc177;
  wire multm_reduce_mulb0_pc178;
  wire multm_reduce_mulb0_pc179;
  wire multm_reduce_mulb0_pc180;
  wire multm_reduce_mulb0_pc181;
  wire multm_reduce_mulb0_pc182;
  wire multm_reduce_mulb0_pc183;
  wire multm_reduce_mulb0_pc184;
  wire multm_reduce_mulb0_ps0;
  wire multm_reduce_mulb0_ps1;
  wire multm_reduce_mulb0_ps2;
  wire multm_reduce_mulb0_ps3;
  wire multm_reduce_mulb0_ps4;
  wire multm_reduce_mulb0_ps5;
  wire multm_reduce_mulb0_ps6;
  wire multm_reduce_mulb0_ps7;
  wire multm_reduce_mulb0_ps8;
  wire multm_reduce_mulb0_ps9;
  wire multm_reduce_mulb0_ps10;
  wire multm_reduce_mulb0_ps11;
  wire multm_reduce_mulb0_ps12;
  wire multm_reduce_mulb0_ps13;
  wire multm_reduce_mulb0_ps14;
  wire multm_reduce_mulb0_ps15;
  wire multm_reduce_mulb0_ps16;
  wire multm_reduce_mulb0_ps17;
  wire multm_reduce_mulb0_ps18;
  wire multm_reduce_mulb0_ps19;
  wire multm_reduce_mulb0_ps20;
  wire multm_reduce_mulb0_ps21;
  wire multm_reduce_mulb0_ps22;
  wire multm_reduce_mulb0_ps23;
  wire multm_reduce_mulb0_ps24;
  wire multm_reduce_mulb0_ps25;
  wire multm_reduce_mulb0_ps26;
  wire multm_reduce_mulb0_ps27;
  wire multm_reduce_mulb0_ps28;
  wire multm_reduce_mulb0_ps29;
  wire multm_reduce_mulb0_ps30;
  wire multm_reduce_mulb0_ps31;
  wire multm_reduce_mulb0_ps32;
  wire multm_reduce_mulb0_ps33;
  wire multm_reduce_mulb0_ps34;
  wire multm_reduce_mulb0_ps35;
  wire multm_reduce_mulb0_ps36;
  wire multm_reduce_mulb0_ps37;
  wire multm_reduce_mulb0_ps38;
  wire multm_reduce_mulb0_ps39;
  wire multm_reduce_mulb0_ps40;
  wire multm_reduce_mulb0_ps41;
  wire multm_reduce_mulb0_ps42;
  wire multm_reduce_mulb0_ps43;
  wire multm_reduce_mulb0_ps44;
  wire multm_reduce_mulb0_ps45;
  wire multm_reduce_mulb0_ps46;
  wire multm_reduce_mulb0_ps47;
  wire multm_reduce_mulb0_ps48;
  wire multm_reduce_mulb0_ps49;
  wire multm_reduce_mulb0_ps50;
  wire multm_reduce_mulb0_ps51;
  wire multm_reduce_mulb0_ps52;
  wire multm_reduce_mulb0_ps53;
  wire multm_reduce_mulb0_ps54;
  wire multm_reduce_mulb0_ps55;
  wire multm_reduce_mulb0_ps56;
  wire multm_reduce_mulb0_ps57;
  wire multm_reduce_mulb0_ps58;
  wire multm_reduce_mulb0_ps59;
  wire multm_reduce_mulb0_ps60;
  wire multm_reduce_mulb0_ps61;
  wire multm_reduce_mulb0_ps62;
  wire multm_reduce_mulb0_ps63;
  wire multm_reduce_mulb0_ps64;
  wire multm_reduce_mulb0_ps65;
  wire multm_reduce_mulb0_ps66;
  wire multm_reduce_mulb0_ps67;
  wire multm_reduce_mulb0_ps68;
  wire multm_reduce_mulb0_ps69;
  wire multm_reduce_mulb0_ps70;
  wire multm_reduce_mulb0_ps71;
  wire multm_reduce_mulb0_ps72;
  wire multm_reduce_mulb0_ps73;
  wire multm_reduce_mulb0_ps74;
  wire multm_reduce_mulb0_ps75;
  wire multm_reduce_mulb0_ps76;
  wire multm_reduce_mulb0_ps77;
  wire multm_reduce_mulb0_ps78;
  wire multm_reduce_mulb0_ps79;
  wire multm_reduce_mulb0_ps80;
  wire multm_reduce_mulb0_ps81;
  wire multm_reduce_mulb0_ps82;
  wire multm_reduce_mulb0_ps83;
  wire multm_reduce_mulb0_ps84;
  wire multm_reduce_mulb0_ps85;
  wire multm_reduce_mulb0_ps86;
  wire multm_reduce_mulb0_ps87;
  wire multm_reduce_mulb0_ps88;
  wire multm_reduce_mulb0_ps89;
  wire multm_reduce_mulb0_ps90;
  wire multm_reduce_mulb0_ps91;
  wire multm_reduce_mulb0_ps92;
  wire multm_reduce_mulb0_ps93;
  wire multm_reduce_mulb0_ps94;
  wire multm_reduce_mulb0_ps95;
  wire multm_reduce_mulb0_ps96;
  wire multm_reduce_mulb0_ps97;
  wire multm_reduce_mulb0_ps98;
  wire multm_reduce_mulb0_ps99;
  wire multm_reduce_mulb0_ps100;
  wire multm_reduce_mulb0_ps101;
  wire multm_reduce_mulb0_ps102;
  wire multm_reduce_mulb0_ps103;
  wire multm_reduce_mulb0_ps104;
  wire multm_reduce_mulb0_ps105;
  wire multm_reduce_mulb0_ps106;
  wire multm_reduce_mulb0_ps107;
  wire multm_reduce_mulb0_ps108;
  wire multm_reduce_mulb0_ps109;
  wire multm_reduce_mulb0_ps110;
  wire multm_reduce_mulb0_ps111;
  wire multm_reduce_mulb0_ps112;
  wire multm_reduce_mulb0_ps113;
  wire multm_reduce_mulb0_ps114;
  wire multm_reduce_mulb0_ps115;
  wire multm_reduce_mulb0_ps116;
  wire multm_reduce_mulb0_ps117;
  wire multm_reduce_mulb0_ps118;
  wire multm_reduce_mulb0_ps119;
  wire multm_reduce_mulb0_ps120;
  wire multm_reduce_mulb0_ps121;
  wire multm_reduce_mulb0_ps122;
  wire multm_reduce_mulb0_ps123;
  wire multm_reduce_mulb0_ps124;
  wire multm_reduce_mulb0_ps125;
  wire multm_reduce_mulb0_ps126;
  wire multm_reduce_mulb0_ps127;
  wire multm_reduce_mulb0_ps128;
  wire multm_reduce_mulb0_ps129;
  wire multm_reduce_mulb0_ps130;
  wire multm_reduce_mulb0_ps131;
  wire multm_reduce_mulb0_ps132;
  wire multm_reduce_mulb0_ps133;
  wire multm_reduce_mulb0_ps134;
  wire multm_reduce_mulb0_ps135;
  wire multm_reduce_mulb0_ps136;
  wire multm_reduce_mulb0_ps137;
  wire multm_reduce_mulb0_ps138;
  wire multm_reduce_mulb0_ps139;
  wire multm_reduce_mulb0_ps140;
  wire multm_reduce_mulb0_ps141;
  wire multm_reduce_mulb0_ps142;
  wire multm_reduce_mulb0_ps143;
  wire multm_reduce_mulb0_ps144;
  wire multm_reduce_mulb0_ps145;
  wire multm_reduce_mulb0_ps146;
  wire multm_reduce_mulb0_ps147;
  wire multm_reduce_mulb0_ps148;
  wire multm_reduce_mulb0_ps149;
  wire multm_reduce_mulb0_ps150;
  wire multm_reduce_mulb0_ps151;
  wire multm_reduce_mulb0_ps152;
  wire multm_reduce_mulb0_ps153;
  wire multm_reduce_mulb0_ps154;
  wire multm_reduce_mulb0_ps155;
  wire multm_reduce_mulb0_ps156;
  wire multm_reduce_mulb0_ps157;
  wire multm_reduce_mulb0_ps158;
  wire multm_reduce_mulb0_ps159;
  wire multm_reduce_mulb0_ps160;
  wire multm_reduce_mulb0_ps161;
  wire multm_reduce_mulb0_ps162;
  wire multm_reduce_mulb0_ps163;
  wire multm_reduce_mulb0_ps164;
  wire multm_reduce_mulb0_ps165;
  wire multm_reduce_mulb0_ps166;
  wire multm_reduce_mulb0_ps167;
  wire multm_reduce_mulb0_ps168;
  wire multm_reduce_mulb0_ps169;
  wire multm_reduce_mulb0_ps170;
  wire multm_reduce_mulb0_ps171;
  wire multm_reduce_mulb0_ps172;
  wire multm_reduce_mulb0_ps173;
  wire multm_reduce_mulb0_ps174;
  wire multm_reduce_mulb0_ps175;
  wire multm_reduce_mulb0_ps176;
  wire multm_reduce_mulb0_ps177;
  wire multm_reduce_mulb0_ps178;
  wire multm_reduce_mulb0_ps179;
  wire multm_reduce_mulb0_ps180;
  wire multm_reduce_mulb0_ps181;
  wire multm_reduce_mulb0_ps182;
  wire multm_reduce_mulb0_ps183;
  wire multm_reduce_mulb0_sq0;
  wire multm_reduce_mulb0_sq1;
  wire multm_reduce_mulb0_sq2;
  wire multm_reduce_mulb0_sq3;
  wire multm_reduce_mulb0_sq4;
  wire multm_reduce_mulb0_sq5;
  wire multm_reduce_mulb0_sq6;
  wire multm_reduce_mulb0_sq7;
  wire multm_reduce_mulb0_sq8;
  wire multm_reduce_mulb0_sq9;
  wire multm_reduce_mulb0_sq10;
  wire multm_reduce_mulb0_sq11;
  wire multm_reduce_mulb0_sq12;
  wire multm_reduce_mulb0_sq13;
  wire multm_reduce_mulb0_sq14;
  wire multm_reduce_mulb0_sq15;
  wire multm_reduce_mulb0_sq16;
  wire multm_reduce_mulb0_sq17;
  wire multm_reduce_mulb0_sq18;
  wire multm_reduce_mulb0_sq19;
  wire multm_reduce_mulb0_sq20;
  wire multm_reduce_mulb0_sq21;
  wire multm_reduce_mulb0_sq22;
  wire multm_reduce_mulb0_sq23;
  wire multm_reduce_mulb0_sq24;
  wire multm_reduce_mulb0_sq25;
  wire multm_reduce_mulb0_sq26;
  wire multm_reduce_mulb0_sq27;
  wire multm_reduce_mulb0_sq28;
  wire multm_reduce_mulb0_sq29;
  wire multm_reduce_mulb0_sq30;
  wire multm_reduce_mulb0_sq31;
  wire multm_reduce_mulb0_sq32;
  wire multm_reduce_mulb0_sq33;
  wire multm_reduce_mulb0_sq34;
  wire multm_reduce_mulb0_sq35;
  wire multm_reduce_mulb0_sq36;
  wire multm_reduce_mulb0_sq37;
  wire multm_reduce_mulb0_sq38;
  wire multm_reduce_mulb0_sq39;
  wire multm_reduce_mulb0_sq40;
  wire multm_reduce_mulb0_sq41;
  wire multm_reduce_mulb0_sq42;
  wire multm_reduce_mulb0_sq43;
  wire multm_reduce_mulb0_sq44;
  wire multm_reduce_mulb0_sq45;
  wire multm_reduce_mulb0_sq46;
  wire multm_reduce_mulb0_sq47;
  wire multm_reduce_mulb0_sq48;
  wire multm_reduce_mulb0_sq49;
  wire multm_reduce_mulb0_sq50;
  wire multm_reduce_mulb0_sq51;
  wire multm_reduce_mulb0_sq52;
  wire multm_reduce_mulb0_sq53;
  wire multm_reduce_mulb0_sq54;
  wire multm_reduce_mulb0_sq55;
  wire multm_reduce_mulb0_sq56;
  wire multm_reduce_mulb0_sq57;
  wire multm_reduce_mulb0_sq58;
  wire multm_reduce_mulb0_sq59;
  wire multm_reduce_mulb0_sq60;
  wire multm_reduce_mulb0_sq61;
  wire multm_reduce_mulb0_sq62;
  wire multm_reduce_mulb0_sq63;
  wire multm_reduce_mulb0_sq64;
  wire multm_reduce_mulb0_sq65;
  wire multm_reduce_mulb0_sq66;
  wire multm_reduce_mulb0_sq67;
  wire multm_reduce_mulb0_sq68;
  wire multm_reduce_mulb0_sq69;
  wire multm_reduce_mulb0_sq70;
  wire multm_reduce_mulb0_sq71;
  wire multm_reduce_mulb0_sq72;
  wire multm_reduce_mulb0_sq73;
  wire multm_reduce_mulb0_sq74;
  wire multm_reduce_mulb0_sq75;
  wire multm_reduce_mulb0_sq76;
  wire multm_reduce_mulb0_sq77;
  wire multm_reduce_mulb0_sq78;
  wire multm_reduce_mulb0_sq79;
  wire multm_reduce_mulb0_sq80;
  wire multm_reduce_mulb0_sq81;
  wire multm_reduce_mulb0_sq82;
  wire multm_reduce_mulb0_sq83;
  wire multm_reduce_mulb0_sq84;
  wire multm_reduce_mulb0_sq85;
  wire multm_reduce_mulb0_sq86;
  wire multm_reduce_mulb0_sq87;
  wire multm_reduce_mulb0_sq88;
  wire multm_reduce_mulb0_sq89;
  wire multm_reduce_mulb0_sq90;
  wire multm_reduce_mulb0_sq91;
  wire multm_reduce_mulb0_sq92;
  wire multm_reduce_mulb0_sq93;
  wire multm_reduce_mulb0_sq94;
  wire multm_reduce_mulb0_sq95;
  wire multm_reduce_mulb0_sq96;
  wire multm_reduce_mulb0_sq97;
  wire multm_reduce_mulb0_sq98;
  wire multm_reduce_mulb0_sq99;
  wire multm_reduce_mulb0_sq100;
  wire multm_reduce_mulb0_sq101;
  wire multm_reduce_mulb0_sq102;
  wire multm_reduce_mulb0_sq103;
  wire multm_reduce_mulb0_sq104;
  wire multm_reduce_mulb0_sq105;
  wire multm_reduce_mulb0_sq106;
  wire multm_reduce_mulb0_sq107;
  wire multm_reduce_mulb0_sq108;
  wire multm_reduce_mulb0_sq109;
  wire multm_reduce_mulb0_sq110;
  wire multm_reduce_mulb0_sq111;
  wire multm_reduce_mulb0_sq112;
  wire multm_reduce_mulb0_sq113;
  wire multm_reduce_mulb0_sq114;
  wire multm_reduce_mulb0_sq115;
  wire multm_reduce_mulb0_sq116;
  wire multm_reduce_mulb0_sq117;
  wire multm_reduce_mulb0_sq118;
  wire multm_reduce_mulb0_sq119;
  wire multm_reduce_mulb0_sq120;
  wire multm_reduce_mulb0_sq121;
  wire multm_reduce_mulb0_sq122;
  wire multm_reduce_mulb0_sq123;
  wire multm_reduce_mulb0_sq124;
  wire multm_reduce_mulb0_sq125;
  wire multm_reduce_mulb0_sq126;
  wire multm_reduce_mulb0_sq127;
  wire multm_reduce_mulb0_sq128;
  wire multm_reduce_mulb0_sq129;
  wire multm_reduce_mulb0_sq130;
  wire multm_reduce_mulb0_sq131;
  wire multm_reduce_mulb0_sq132;
  wire multm_reduce_mulb0_sq133;
  wire multm_reduce_mulb0_sq134;
  wire multm_reduce_mulb0_sq135;
  wire multm_reduce_mulb0_sq136;
  wire multm_reduce_mulb0_sq137;
  wire multm_reduce_mulb0_sq138;
  wire multm_reduce_mulb0_sq139;
  wire multm_reduce_mulb0_sq140;
  wire multm_reduce_mulb0_sq141;
  wire multm_reduce_mulb0_sq142;
  wire multm_reduce_mulb0_sq143;
  wire multm_reduce_mulb0_sq144;
  wire multm_reduce_mulb0_sq145;
  wire multm_reduce_mulb0_sq146;
  wire multm_reduce_mulb0_sq147;
  wire multm_reduce_mulb0_sq148;
  wire multm_reduce_mulb0_sq149;
  wire multm_reduce_mulb0_sq150;
  wire multm_reduce_mulb0_sq151;
  wire multm_reduce_mulb0_sq152;
  wire multm_reduce_mulb0_sq153;
  wire multm_reduce_mulb0_sq154;
  wire multm_reduce_mulb0_sq155;
  wire multm_reduce_mulb0_sq156;
  wire multm_reduce_mulb0_sq157;
  wire multm_reduce_mulb0_sq158;
  wire multm_reduce_mulb0_sq159;
  wire multm_reduce_mulb0_sq160;
  wire multm_reduce_mulb0_sq161;
  wire multm_reduce_mulb0_sq162;
  wire multm_reduce_mulb0_sq163;
  wire multm_reduce_mulb0_sq164;
  wire multm_reduce_mulb0_sq165;
  wire multm_reduce_mulb0_sq166;
  wire multm_reduce_mulb0_sq167;
  wire multm_reduce_mulb0_sq168;
  wire multm_reduce_mulb0_sq169;
  wire multm_reduce_mulb0_sq170;
  wire multm_reduce_mulb0_sq171;
  wire multm_reduce_mulb0_sq172;
  wire multm_reduce_mulb0_sq173;
  wire multm_reduce_mulb0_sq174;
  wire multm_reduce_mulb0_sq175;
  wire multm_reduce_mulb0_sq176;
  wire multm_reduce_mulb0_sq177;
  wire multm_reduce_mulb0_sq178;
  wire multm_reduce_mulb0_sq179;
  wire multm_reduce_mulb0_sq180;
  wire multm_reduce_mulb0_sq181;
  wire multm_reduce_mulb0_sq182;
  wire multm_reduce_mulb0_sq183;
  wire multm_reduce_mulb0_sq184;
  wire multm_reduce_mulb1_add3_maj3_or3_wx;
  wire multm_reduce_mulb1_add3_maj3_wx;
  wire multm_reduce_mulb1_add3_maj3_wy;
  wire multm_reduce_mulb1_add3_maj3_xy;
  wire multm_reduce_mulb1_add3_xor3_wx;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx0;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx1;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx4;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx5;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx6;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx7;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx10;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx12;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx18;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx20;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx22;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx23;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx24;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx28;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx30;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx32;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx34;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx37;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx40;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx41;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx42;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx43;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx47;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx48;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx51;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx52;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx53;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx54;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx55;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx57;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx62;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx66;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx68;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx69;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx71;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx73;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx74;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx79;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx80;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx82;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx86;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx88;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx90;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx91;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx96;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx99;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx100;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx101;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx102;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx104;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx105;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx107;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx108;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx109;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx110;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx112;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx114;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx117;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx118;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx119;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx120;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx121;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx122;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx123;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx128;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx130;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx132;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx135;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx136;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx140;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx141;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx142;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx143;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx144;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx147;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx150;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx151;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx152;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx153;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx155;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx156;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx157;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx158;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx159;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx160;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx162;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx166;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx171;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx172;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx173;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx174;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx175;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx179;
  wire multm_reduce_mulb1_add3b_maj3b_or3b_wx181;
  wire multm_reduce_mulb1_add3b_maj3b_wx0;
  wire multm_reduce_mulb1_add3b_maj3b_wx1;
  wire multm_reduce_mulb1_add3b_maj3b_wx4;
  wire multm_reduce_mulb1_add3b_maj3b_wx5;
  wire multm_reduce_mulb1_add3b_maj3b_wx6;
  wire multm_reduce_mulb1_add3b_maj3b_wx7;
  wire multm_reduce_mulb1_add3b_maj3b_wx10;
  wire multm_reduce_mulb1_add3b_maj3b_wx12;
  wire multm_reduce_mulb1_add3b_maj3b_wx18;
  wire multm_reduce_mulb1_add3b_maj3b_wx20;
  wire multm_reduce_mulb1_add3b_maj3b_wx22;
  wire multm_reduce_mulb1_add3b_maj3b_wx23;
  wire multm_reduce_mulb1_add3b_maj3b_wx24;
  wire multm_reduce_mulb1_add3b_maj3b_wx28;
  wire multm_reduce_mulb1_add3b_maj3b_wx30;
  wire multm_reduce_mulb1_add3b_maj3b_wx32;
  wire multm_reduce_mulb1_add3b_maj3b_wx34;
  wire multm_reduce_mulb1_add3b_maj3b_wx37;
  wire multm_reduce_mulb1_add3b_maj3b_wx40;
  wire multm_reduce_mulb1_add3b_maj3b_wx41;
  wire multm_reduce_mulb1_add3b_maj3b_wx42;
  wire multm_reduce_mulb1_add3b_maj3b_wx43;
  wire multm_reduce_mulb1_add3b_maj3b_wx47;
  wire multm_reduce_mulb1_add3b_maj3b_wx48;
  wire multm_reduce_mulb1_add3b_maj3b_wx51;
  wire multm_reduce_mulb1_add3b_maj3b_wx52;
  wire multm_reduce_mulb1_add3b_maj3b_wx53;
  wire multm_reduce_mulb1_add3b_maj3b_wx54;
  wire multm_reduce_mulb1_add3b_maj3b_wx55;
  wire multm_reduce_mulb1_add3b_maj3b_wx57;
  wire multm_reduce_mulb1_add3b_maj3b_wx62;
  wire multm_reduce_mulb1_add3b_maj3b_wx66;
  wire multm_reduce_mulb1_add3b_maj3b_wx68;
  wire multm_reduce_mulb1_add3b_maj3b_wx69;
  wire multm_reduce_mulb1_add3b_maj3b_wx71;
  wire multm_reduce_mulb1_add3b_maj3b_wx73;
  wire multm_reduce_mulb1_add3b_maj3b_wx74;
  wire multm_reduce_mulb1_add3b_maj3b_wx79;
  wire multm_reduce_mulb1_add3b_maj3b_wx80;
  wire multm_reduce_mulb1_add3b_maj3b_wx82;
  wire multm_reduce_mulb1_add3b_maj3b_wx86;
  wire multm_reduce_mulb1_add3b_maj3b_wx88;
  wire multm_reduce_mulb1_add3b_maj3b_wx90;
  wire multm_reduce_mulb1_add3b_maj3b_wx91;
  wire multm_reduce_mulb1_add3b_maj3b_wx96;
  wire multm_reduce_mulb1_add3b_maj3b_wx99;
  wire multm_reduce_mulb1_add3b_maj3b_wx100;
  wire multm_reduce_mulb1_add3b_maj3b_wx101;
  wire multm_reduce_mulb1_add3b_maj3b_wx102;
  wire multm_reduce_mulb1_add3b_maj3b_wx104;
  wire multm_reduce_mulb1_add3b_maj3b_wx105;
  wire multm_reduce_mulb1_add3b_maj3b_wx107;
  wire multm_reduce_mulb1_add3b_maj3b_wx108;
  wire multm_reduce_mulb1_add3b_maj3b_wx109;
  wire multm_reduce_mulb1_add3b_maj3b_wx110;
  wire multm_reduce_mulb1_add3b_maj3b_wx112;
  wire multm_reduce_mulb1_add3b_maj3b_wx114;
  wire multm_reduce_mulb1_add3b_maj3b_wx117;
  wire multm_reduce_mulb1_add3b_maj3b_wx118;
  wire multm_reduce_mulb1_add3b_maj3b_wx119;
  wire multm_reduce_mulb1_add3b_maj3b_wx120;
  wire multm_reduce_mulb1_add3b_maj3b_wx121;
  wire multm_reduce_mulb1_add3b_maj3b_wx122;
  wire multm_reduce_mulb1_add3b_maj3b_wx123;
  wire multm_reduce_mulb1_add3b_maj3b_wx128;
  wire multm_reduce_mulb1_add3b_maj3b_wx130;
  wire multm_reduce_mulb1_add3b_maj3b_wx132;
  wire multm_reduce_mulb1_add3b_maj3b_wx135;
  wire multm_reduce_mulb1_add3b_maj3b_wx136;
  wire multm_reduce_mulb1_add3b_maj3b_wx140;
  wire multm_reduce_mulb1_add3b_maj3b_wx141;
  wire multm_reduce_mulb1_add3b_maj3b_wx142;
  wire multm_reduce_mulb1_add3b_maj3b_wx143;
  wire multm_reduce_mulb1_add3b_maj3b_wx144;
  wire multm_reduce_mulb1_add3b_maj3b_wx147;
  wire multm_reduce_mulb1_add3b_maj3b_wx150;
  wire multm_reduce_mulb1_add3b_maj3b_wx151;
  wire multm_reduce_mulb1_add3b_maj3b_wx152;
  wire multm_reduce_mulb1_add3b_maj3b_wx153;
  wire multm_reduce_mulb1_add3b_maj3b_wx155;
  wire multm_reduce_mulb1_add3b_maj3b_wx156;
  wire multm_reduce_mulb1_add3b_maj3b_wx157;
  wire multm_reduce_mulb1_add3b_maj3b_wx158;
  wire multm_reduce_mulb1_add3b_maj3b_wx159;
  wire multm_reduce_mulb1_add3b_maj3b_wx160;
  wire multm_reduce_mulb1_add3b_maj3b_wx162;
  wire multm_reduce_mulb1_add3b_maj3b_wx166;
  wire multm_reduce_mulb1_add3b_maj3b_wx171;
  wire multm_reduce_mulb1_add3b_maj3b_wx172;
  wire multm_reduce_mulb1_add3b_maj3b_wx173;
  wire multm_reduce_mulb1_add3b_maj3b_wx174;
  wire multm_reduce_mulb1_add3b_maj3b_wx175;
  wire multm_reduce_mulb1_add3b_maj3b_wx179;
  wire multm_reduce_mulb1_add3b_maj3b_wx181;
  wire multm_reduce_mulb1_add3b_maj3b_wy0;
  wire multm_reduce_mulb1_add3b_maj3b_wy1;
  wire multm_reduce_mulb1_add3b_maj3b_wy4;
  wire multm_reduce_mulb1_add3b_maj3b_wy5;
  wire multm_reduce_mulb1_add3b_maj3b_wy6;
  wire multm_reduce_mulb1_add3b_maj3b_wy7;
  wire multm_reduce_mulb1_add3b_maj3b_wy10;
  wire multm_reduce_mulb1_add3b_maj3b_wy12;
  wire multm_reduce_mulb1_add3b_maj3b_wy18;
  wire multm_reduce_mulb1_add3b_maj3b_wy20;
  wire multm_reduce_mulb1_add3b_maj3b_wy22;
  wire multm_reduce_mulb1_add3b_maj3b_wy23;
  wire multm_reduce_mulb1_add3b_maj3b_wy24;
  wire multm_reduce_mulb1_add3b_maj3b_wy28;
  wire multm_reduce_mulb1_add3b_maj3b_wy30;
  wire multm_reduce_mulb1_add3b_maj3b_wy32;
  wire multm_reduce_mulb1_add3b_maj3b_wy34;
  wire multm_reduce_mulb1_add3b_maj3b_wy37;
  wire multm_reduce_mulb1_add3b_maj3b_wy40;
  wire multm_reduce_mulb1_add3b_maj3b_wy41;
  wire multm_reduce_mulb1_add3b_maj3b_wy42;
  wire multm_reduce_mulb1_add3b_maj3b_wy43;
  wire multm_reduce_mulb1_add3b_maj3b_wy47;
  wire multm_reduce_mulb1_add3b_maj3b_wy48;
  wire multm_reduce_mulb1_add3b_maj3b_wy51;
  wire multm_reduce_mulb1_add3b_maj3b_wy52;
  wire multm_reduce_mulb1_add3b_maj3b_wy53;
  wire multm_reduce_mulb1_add3b_maj3b_wy54;
  wire multm_reduce_mulb1_add3b_maj3b_wy55;
  wire multm_reduce_mulb1_add3b_maj3b_wy57;
  wire multm_reduce_mulb1_add3b_maj3b_wy62;
  wire multm_reduce_mulb1_add3b_maj3b_wy66;
  wire multm_reduce_mulb1_add3b_maj3b_wy68;
  wire multm_reduce_mulb1_add3b_maj3b_wy69;
  wire multm_reduce_mulb1_add3b_maj3b_wy71;
  wire multm_reduce_mulb1_add3b_maj3b_wy73;
  wire multm_reduce_mulb1_add3b_maj3b_wy74;
  wire multm_reduce_mulb1_add3b_maj3b_wy79;
  wire multm_reduce_mulb1_add3b_maj3b_wy80;
  wire multm_reduce_mulb1_add3b_maj3b_wy82;
  wire multm_reduce_mulb1_add3b_maj3b_wy86;
  wire multm_reduce_mulb1_add3b_maj3b_wy88;
  wire multm_reduce_mulb1_add3b_maj3b_wy90;
  wire multm_reduce_mulb1_add3b_maj3b_wy91;
  wire multm_reduce_mulb1_add3b_maj3b_wy96;
  wire multm_reduce_mulb1_add3b_maj3b_wy99;
  wire multm_reduce_mulb1_add3b_maj3b_wy100;
  wire multm_reduce_mulb1_add3b_maj3b_wy101;
  wire multm_reduce_mulb1_add3b_maj3b_wy102;
  wire multm_reduce_mulb1_add3b_maj3b_wy104;
  wire multm_reduce_mulb1_add3b_maj3b_wy105;
  wire multm_reduce_mulb1_add3b_maj3b_wy107;
  wire multm_reduce_mulb1_add3b_maj3b_wy108;
  wire multm_reduce_mulb1_add3b_maj3b_wy109;
  wire multm_reduce_mulb1_add3b_maj3b_wy110;
  wire multm_reduce_mulb1_add3b_maj3b_wy112;
  wire multm_reduce_mulb1_add3b_maj3b_wy114;
  wire multm_reduce_mulb1_add3b_maj3b_wy117;
  wire multm_reduce_mulb1_add3b_maj3b_wy118;
  wire multm_reduce_mulb1_add3b_maj3b_wy119;
  wire multm_reduce_mulb1_add3b_maj3b_wy120;
  wire multm_reduce_mulb1_add3b_maj3b_wy121;
  wire multm_reduce_mulb1_add3b_maj3b_wy122;
  wire multm_reduce_mulb1_add3b_maj3b_wy123;
  wire multm_reduce_mulb1_add3b_maj3b_wy128;
  wire multm_reduce_mulb1_add3b_maj3b_wy130;
  wire multm_reduce_mulb1_add3b_maj3b_wy132;
  wire multm_reduce_mulb1_add3b_maj3b_wy135;
  wire multm_reduce_mulb1_add3b_maj3b_wy136;
  wire multm_reduce_mulb1_add3b_maj3b_wy140;
  wire multm_reduce_mulb1_add3b_maj3b_wy141;
  wire multm_reduce_mulb1_add3b_maj3b_wy142;
  wire multm_reduce_mulb1_add3b_maj3b_wy143;
  wire multm_reduce_mulb1_add3b_maj3b_wy144;
  wire multm_reduce_mulb1_add3b_maj3b_wy147;
  wire multm_reduce_mulb1_add3b_maj3b_wy150;
  wire multm_reduce_mulb1_add3b_maj3b_wy151;
  wire multm_reduce_mulb1_add3b_maj3b_wy152;
  wire multm_reduce_mulb1_add3b_maj3b_wy153;
  wire multm_reduce_mulb1_add3b_maj3b_wy155;
  wire multm_reduce_mulb1_add3b_maj3b_wy156;
  wire multm_reduce_mulb1_add3b_maj3b_wy157;
  wire multm_reduce_mulb1_add3b_maj3b_wy158;
  wire multm_reduce_mulb1_add3b_maj3b_wy159;
  wire multm_reduce_mulb1_add3b_maj3b_wy160;
  wire multm_reduce_mulb1_add3b_maj3b_wy162;
  wire multm_reduce_mulb1_add3b_maj3b_wy166;
  wire multm_reduce_mulb1_add3b_maj3b_wy171;
  wire multm_reduce_mulb1_add3b_maj3b_wy172;
  wire multm_reduce_mulb1_add3b_maj3b_wy173;
  wire multm_reduce_mulb1_add3b_maj3b_wy174;
  wire multm_reduce_mulb1_add3b_maj3b_wy175;
  wire multm_reduce_mulb1_add3b_maj3b_wy179;
  wire multm_reduce_mulb1_add3b_maj3b_wy181;
  wire multm_reduce_mulb1_add3b_maj3b_xy0;
  wire multm_reduce_mulb1_add3b_maj3b_xy1;
  wire multm_reduce_mulb1_add3b_maj3b_xy4;
  wire multm_reduce_mulb1_add3b_maj3b_xy5;
  wire multm_reduce_mulb1_add3b_maj3b_xy6;
  wire multm_reduce_mulb1_add3b_maj3b_xy7;
  wire multm_reduce_mulb1_add3b_maj3b_xy10;
  wire multm_reduce_mulb1_add3b_maj3b_xy12;
  wire multm_reduce_mulb1_add3b_maj3b_xy18;
  wire multm_reduce_mulb1_add3b_maj3b_xy20;
  wire multm_reduce_mulb1_add3b_maj3b_xy22;
  wire multm_reduce_mulb1_add3b_maj3b_xy23;
  wire multm_reduce_mulb1_add3b_maj3b_xy24;
  wire multm_reduce_mulb1_add3b_maj3b_xy28;
  wire multm_reduce_mulb1_add3b_maj3b_xy30;
  wire multm_reduce_mulb1_add3b_maj3b_xy32;
  wire multm_reduce_mulb1_add3b_maj3b_xy34;
  wire multm_reduce_mulb1_add3b_maj3b_xy37;
  wire multm_reduce_mulb1_add3b_maj3b_xy40;
  wire multm_reduce_mulb1_add3b_maj3b_xy41;
  wire multm_reduce_mulb1_add3b_maj3b_xy42;
  wire multm_reduce_mulb1_add3b_maj3b_xy43;
  wire multm_reduce_mulb1_add3b_maj3b_xy47;
  wire multm_reduce_mulb1_add3b_maj3b_xy48;
  wire multm_reduce_mulb1_add3b_maj3b_xy51;
  wire multm_reduce_mulb1_add3b_maj3b_xy52;
  wire multm_reduce_mulb1_add3b_maj3b_xy53;
  wire multm_reduce_mulb1_add3b_maj3b_xy54;
  wire multm_reduce_mulb1_add3b_maj3b_xy55;
  wire multm_reduce_mulb1_add3b_maj3b_xy57;
  wire multm_reduce_mulb1_add3b_maj3b_xy62;
  wire multm_reduce_mulb1_add3b_maj3b_xy66;
  wire multm_reduce_mulb1_add3b_maj3b_xy68;
  wire multm_reduce_mulb1_add3b_maj3b_xy69;
  wire multm_reduce_mulb1_add3b_maj3b_xy71;
  wire multm_reduce_mulb1_add3b_maj3b_xy73;
  wire multm_reduce_mulb1_add3b_maj3b_xy74;
  wire multm_reduce_mulb1_add3b_maj3b_xy79;
  wire multm_reduce_mulb1_add3b_maj3b_xy80;
  wire multm_reduce_mulb1_add3b_maj3b_xy82;
  wire multm_reduce_mulb1_add3b_maj3b_xy86;
  wire multm_reduce_mulb1_add3b_maj3b_xy88;
  wire multm_reduce_mulb1_add3b_maj3b_xy90;
  wire multm_reduce_mulb1_add3b_maj3b_xy91;
  wire multm_reduce_mulb1_add3b_maj3b_xy96;
  wire multm_reduce_mulb1_add3b_maj3b_xy99;
  wire multm_reduce_mulb1_add3b_maj3b_xy100;
  wire multm_reduce_mulb1_add3b_maj3b_xy101;
  wire multm_reduce_mulb1_add3b_maj3b_xy102;
  wire multm_reduce_mulb1_add3b_maj3b_xy104;
  wire multm_reduce_mulb1_add3b_maj3b_xy105;
  wire multm_reduce_mulb1_add3b_maj3b_xy107;
  wire multm_reduce_mulb1_add3b_maj3b_xy108;
  wire multm_reduce_mulb1_add3b_maj3b_xy109;
  wire multm_reduce_mulb1_add3b_maj3b_xy110;
  wire multm_reduce_mulb1_add3b_maj3b_xy112;
  wire multm_reduce_mulb1_add3b_maj3b_xy114;
  wire multm_reduce_mulb1_add3b_maj3b_xy117;
  wire multm_reduce_mulb1_add3b_maj3b_xy118;
  wire multm_reduce_mulb1_add3b_maj3b_xy119;
  wire multm_reduce_mulb1_add3b_maj3b_xy120;
  wire multm_reduce_mulb1_add3b_maj3b_xy121;
  wire multm_reduce_mulb1_add3b_maj3b_xy122;
  wire multm_reduce_mulb1_add3b_maj3b_xy123;
  wire multm_reduce_mulb1_add3b_maj3b_xy128;
  wire multm_reduce_mulb1_add3b_maj3b_xy130;
  wire multm_reduce_mulb1_add3b_maj3b_xy132;
  wire multm_reduce_mulb1_add3b_maj3b_xy135;
  wire multm_reduce_mulb1_add3b_maj3b_xy136;
  wire multm_reduce_mulb1_add3b_maj3b_xy140;
  wire multm_reduce_mulb1_add3b_maj3b_xy141;
  wire multm_reduce_mulb1_add3b_maj3b_xy142;
  wire multm_reduce_mulb1_add3b_maj3b_xy143;
  wire multm_reduce_mulb1_add3b_maj3b_xy144;
  wire multm_reduce_mulb1_add3b_maj3b_xy147;
  wire multm_reduce_mulb1_add3b_maj3b_xy150;
  wire multm_reduce_mulb1_add3b_maj3b_xy151;
  wire multm_reduce_mulb1_add3b_maj3b_xy152;
  wire multm_reduce_mulb1_add3b_maj3b_xy153;
  wire multm_reduce_mulb1_add3b_maj3b_xy155;
  wire multm_reduce_mulb1_add3b_maj3b_xy156;
  wire multm_reduce_mulb1_add3b_maj3b_xy157;
  wire multm_reduce_mulb1_add3b_maj3b_xy158;
  wire multm_reduce_mulb1_add3b_maj3b_xy159;
  wire multm_reduce_mulb1_add3b_maj3b_xy160;
  wire multm_reduce_mulb1_add3b_maj3b_xy162;
  wire multm_reduce_mulb1_add3b_maj3b_xy166;
  wire multm_reduce_mulb1_add3b_maj3b_xy171;
  wire multm_reduce_mulb1_add3b_maj3b_xy172;
  wire multm_reduce_mulb1_add3b_maj3b_xy173;
  wire multm_reduce_mulb1_add3b_maj3b_xy174;
  wire multm_reduce_mulb1_add3b_maj3b_xy175;
  wire multm_reduce_mulb1_add3b_maj3b_xy179;
  wire multm_reduce_mulb1_add3b_maj3b_xy181;
  wire multm_reduce_mulb1_add3b_xor3b_wx0;
  wire multm_reduce_mulb1_add3b_xor3b_wx1;
  wire multm_reduce_mulb1_add3b_xor3b_wx4;
  wire multm_reduce_mulb1_add3b_xor3b_wx5;
  wire multm_reduce_mulb1_add3b_xor3b_wx6;
  wire multm_reduce_mulb1_add3b_xor3b_wx7;
  wire multm_reduce_mulb1_add3b_xor3b_wx10;
  wire multm_reduce_mulb1_add3b_xor3b_wx12;
  wire multm_reduce_mulb1_add3b_xor3b_wx18;
  wire multm_reduce_mulb1_add3b_xor3b_wx20;
  wire multm_reduce_mulb1_add3b_xor3b_wx22;
  wire multm_reduce_mulb1_add3b_xor3b_wx23;
  wire multm_reduce_mulb1_add3b_xor3b_wx24;
  wire multm_reduce_mulb1_add3b_xor3b_wx28;
  wire multm_reduce_mulb1_add3b_xor3b_wx30;
  wire multm_reduce_mulb1_add3b_xor3b_wx32;
  wire multm_reduce_mulb1_add3b_xor3b_wx34;
  wire multm_reduce_mulb1_add3b_xor3b_wx37;
  wire multm_reduce_mulb1_add3b_xor3b_wx40;
  wire multm_reduce_mulb1_add3b_xor3b_wx41;
  wire multm_reduce_mulb1_add3b_xor3b_wx42;
  wire multm_reduce_mulb1_add3b_xor3b_wx43;
  wire multm_reduce_mulb1_add3b_xor3b_wx47;
  wire multm_reduce_mulb1_add3b_xor3b_wx48;
  wire multm_reduce_mulb1_add3b_xor3b_wx51;
  wire multm_reduce_mulb1_add3b_xor3b_wx52;
  wire multm_reduce_mulb1_add3b_xor3b_wx53;
  wire multm_reduce_mulb1_add3b_xor3b_wx54;
  wire multm_reduce_mulb1_add3b_xor3b_wx55;
  wire multm_reduce_mulb1_add3b_xor3b_wx57;
  wire multm_reduce_mulb1_add3b_xor3b_wx62;
  wire multm_reduce_mulb1_add3b_xor3b_wx66;
  wire multm_reduce_mulb1_add3b_xor3b_wx68;
  wire multm_reduce_mulb1_add3b_xor3b_wx69;
  wire multm_reduce_mulb1_add3b_xor3b_wx71;
  wire multm_reduce_mulb1_add3b_xor3b_wx73;
  wire multm_reduce_mulb1_add3b_xor3b_wx74;
  wire multm_reduce_mulb1_add3b_xor3b_wx79;
  wire multm_reduce_mulb1_add3b_xor3b_wx80;
  wire multm_reduce_mulb1_add3b_xor3b_wx82;
  wire multm_reduce_mulb1_add3b_xor3b_wx86;
  wire multm_reduce_mulb1_add3b_xor3b_wx88;
  wire multm_reduce_mulb1_add3b_xor3b_wx90;
  wire multm_reduce_mulb1_add3b_xor3b_wx91;
  wire multm_reduce_mulb1_add3b_xor3b_wx96;
  wire multm_reduce_mulb1_add3b_xor3b_wx99;
  wire multm_reduce_mulb1_add3b_xor3b_wx100;
  wire multm_reduce_mulb1_add3b_xor3b_wx101;
  wire multm_reduce_mulb1_add3b_xor3b_wx102;
  wire multm_reduce_mulb1_add3b_xor3b_wx104;
  wire multm_reduce_mulb1_add3b_xor3b_wx105;
  wire multm_reduce_mulb1_add3b_xor3b_wx107;
  wire multm_reduce_mulb1_add3b_xor3b_wx108;
  wire multm_reduce_mulb1_add3b_xor3b_wx109;
  wire multm_reduce_mulb1_add3b_xor3b_wx110;
  wire multm_reduce_mulb1_add3b_xor3b_wx112;
  wire multm_reduce_mulb1_add3b_xor3b_wx114;
  wire multm_reduce_mulb1_add3b_xor3b_wx117;
  wire multm_reduce_mulb1_add3b_xor3b_wx118;
  wire multm_reduce_mulb1_add3b_xor3b_wx119;
  wire multm_reduce_mulb1_add3b_xor3b_wx120;
  wire multm_reduce_mulb1_add3b_xor3b_wx121;
  wire multm_reduce_mulb1_add3b_xor3b_wx122;
  wire multm_reduce_mulb1_add3b_xor3b_wx123;
  wire multm_reduce_mulb1_add3b_xor3b_wx128;
  wire multm_reduce_mulb1_add3b_xor3b_wx130;
  wire multm_reduce_mulb1_add3b_xor3b_wx132;
  wire multm_reduce_mulb1_add3b_xor3b_wx135;
  wire multm_reduce_mulb1_add3b_xor3b_wx136;
  wire multm_reduce_mulb1_add3b_xor3b_wx140;
  wire multm_reduce_mulb1_add3b_xor3b_wx141;
  wire multm_reduce_mulb1_add3b_xor3b_wx142;
  wire multm_reduce_mulb1_add3b_xor3b_wx143;
  wire multm_reduce_mulb1_add3b_xor3b_wx144;
  wire multm_reduce_mulb1_add3b_xor3b_wx147;
  wire multm_reduce_mulb1_add3b_xor3b_wx150;
  wire multm_reduce_mulb1_add3b_xor3b_wx151;
  wire multm_reduce_mulb1_add3b_xor3b_wx152;
  wire multm_reduce_mulb1_add3b_xor3b_wx153;
  wire multm_reduce_mulb1_add3b_xor3b_wx155;
  wire multm_reduce_mulb1_add3b_xor3b_wx156;
  wire multm_reduce_mulb1_add3b_xor3b_wx157;
  wire multm_reduce_mulb1_add3b_xor3b_wx158;
  wire multm_reduce_mulb1_add3b_xor3b_wx159;
  wire multm_reduce_mulb1_add3b_xor3b_wx160;
  wire multm_reduce_mulb1_add3b_xor3b_wx162;
  wire multm_reduce_mulb1_add3b_xor3b_wx166;
  wire multm_reduce_mulb1_add3b_xor3b_wx171;
  wire multm_reduce_mulb1_add3b_xor3b_wx172;
  wire multm_reduce_mulb1_add3b_xor3b_wx173;
  wire multm_reduce_mulb1_add3b_xor3b_wx174;
  wire multm_reduce_mulb1_add3b_xor3b_wx175;
  wire multm_reduce_mulb1_add3b_xor3b_wx179;
  wire multm_reduce_mulb1_add3b_xor3b_wx181;
  wire multm_reduce_mulb1_cq0;
  wire multm_reduce_mulb1_cq1;
  wire multm_reduce_mulb1_cq2;
  wire multm_reduce_mulb1_cq3;
  wire multm_reduce_mulb1_cq4;
  wire multm_reduce_mulb1_cq5;
  wire multm_reduce_mulb1_cq6;
  wire multm_reduce_mulb1_cq7;
  wire multm_reduce_mulb1_cq8;
  wire multm_reduce_mulb1_cq9;
  wire multm_reduce_mulb1_cq10;
  wire multm_reduce_mulb1_cq11;
  wire multm_reduce_mulb1_cq12;
  wire multm_reduce_mulb1_cq13;
  wire multm_reduce_mulb1_cq14;
  wire multm_reduce_mulb1_cq15;
  wire multm_reduce_mulb1_cq16;
  wire multm_reduce_mulb1_cq17;
  wire multm_reduce_mulb1_cq18;
  wire multm_reduce_mulb1_cq19;
  wire multm_reduce_mulb1_cq20;
  wire multm_reduce_mulb1_cq21;
  wire multm_reduce_mulb1_cq22;
  wire multm_reduce_mulb1_cq23;
  wire multm_reduce_mulb1_cq24;
  wire multm_reduce_mulb1_cq25;
  wire multm_reduce_mulb1_cq26;
  wire multm_reduce_mulb1_cq27;
  wire multm_reduce_mulb1_cq28;
  wire multm_reduce_mulb1_cq29;
  wire multm_reduce_mulb1_cq30;
  wire multm_reduce_mulb1_cq31;
  wire multm_reduce_mulb1_cq32;
  wire multm_reduce_mulb1_cq33;
  wire multm_reduce_mulb1_cq34;
  wire multm_reduce_mulb1_cq35;
  wire multm_reduce_mulb1_cq36;
  wire multm_reduce_mulb1_cq37;
  wire multm_reduce_mulb1_cq38;
  wire multm_reduce_mulb1_cq39;
  wire multm_reduce_mulb1_cq40;
  wire multm_reduce_mulb1_cq41;
  wire multm_reduce_mulb1_cq42;
  wire multm_reduce_mulb1_cq43;
  wire multm_reduce_mulb1_cq44;
  wire multm_reduce_mulb1_cq45;
  wire multm_reduce_mulb1_cq46;
  wire multm_reduce_mulb1_cq47;
  wire multm_reduce_mulb1_cq48;
  wire multm_reduce_mulb1_cq49;
  wire multm_reduce_mulb1_cq50;
  wire multm_reduce_mulb1_cq51;
  wire multm_reduce_mulb1_cq52;
  wire multm_reduce_mulb1_cq53;
  wire multm_reduce_mulb1_cq54;
  wire multm_reduce_mulb1_cq55;
  wire multm_reduce_mulb1_cq56;
  wire multm_reduce_mulb1_cq57;
  wire multm_reduce_mulb1_cq58;
  wire multm_reduce_mulb1_cq59;
  wire multm_reduce_mulb1_cq60;
  wire multm_reduce_mulb1_cq61;
  wire multm_reduce_mulb1_cq62;
  wire multm_reduce_mulb1_cq63;
  wire multm_reduce_mulb1_cq64;
  wire multm_reduce_mulb1_cq65;
  wire multm_reduce_mulb1_cq66;
  wire multm_reduce_mulb1_cq67;
  wire multm_reduce_mulb1_cq68;
  wire multm_reduce_mulb1_cq69;
  wire multm_reduce_mulb1_cq70;
  wire multm_reduce_mulb1_cq71;
  wire multm_reduce_mulb1_cq72;
  wire multm_reduce_mulb1_cq73;
  wire multm_reduce_mulb1_cq74;
  wire multm_reduce_mulb1_cq75;
  wire multm_reduce_mulb1_cq76;
  wire multm_reduce_mulb1_cq77;
  wire multm_reduce_mulb1_cq78;
  wire multm_reduce_mulb1_cq79;
  wire multm_reduce_mulb1_cq80;
  wire multm_reduce_mulb1_cq81;
  wire multm_reduce_mulb1_cq82;
  wire multm_reduce_mulb1_cq83;
  wire multm_reduce_mulb1_cq84;
  wire multm_reduce_mulb1_cq85;
  wire multm_reduce_mulb1_cq86;
  wire multm_reduce_mulb1_cq87;
  wire multm_reduce_mulb1_cq88;
  wire multm_reduce_mulb1_cq89;
  wire multm_reduce_mulb1_cq90;
  wire multm_reduce_mulb1_cq91;
  wire multm_reduce_mulb1_cq92;
  wire multm_reduce_mulb1_cq93;
  wire multm_reduce_mulb1_cq94;
  wire multm_reduce_mulb1_cq95;
  wire multm_reduce_mulb1_cq96;
  wire multm_reduce_mulb1_cq97;
  wire multm_reduce_mulb1_cq98;
  wire multm_reduce_mulb1_cq99;
  wire multm_reduce_mulb1_cq100;
  wire multm_reduce_mulb1_cq101;
  wire multm_reduce_mulb1_cq102;
  wire multm_reduce_mulb1_cq103;
  wire multm_reduce_mulb1_cq104;
  wire multm_reduce_mulb1_cq105;
  wire multm_reduce_mulb1_cq106;
  wire multm_reduce_mulb1_cq107;
  wire multm_reduce_mulb1_cq108;
  wire multm_reduce_mulb1_cq109;
  wire multm_reduce_mulb1_cq110;
  wire multm_reduce_mulb1_cq111;
  wire multm_reduce_mulb1_cq112;
  wire multm_reduce_mulb1_cq113;
  wire multm_reduce_mulb1_cq114;
  wire multm_reduce_mulb1_cq115;
  wire multm_reduce_mulb1_cq116;
  wire multm_reduce_mulb1_cq117;
  wire multm_reduce_mulb1_cq118;
  wire multm_reduce_mulb1_cq119;
  wire multm_reduce_mulb1_cq120;
  wire multm_reduce_mulb1_cq121;
  wire multm_reduce_mulb1_cq122;
  wire multm_reduce_mulb1_cq123;
  wire multm_reduce_mulb1_cq124;
  wire multm_reduce_mulb1_cq125;
  wire multm_reduce_mulb1_cq126;
  wire multm_reduce_mulb1_cq127;
  wire multm_reduce_mulb1_cq128;
  wire multm_reduce_mulb1_cq129;
  wire multm_reduce_mulb1_cq130;
  wire multm_reduce_mulb1_cq131;
  wire multm_reduce_mulb1_cq132;
  wire multm_reduce_mulb1_cq133;
  wire multm_reduce_mulb1_cq134;
  wire multm_reduce_mulb1_cq135;
  wire multm_reduce_mulb1_cq136;
  wire multm_reduce_mulb1_cq137;
  wire multm_reduce_mulb1_cq138;
  wire multm_reduce_mulb1_cq139;
  wire multm_reduce_mulb1_cq140;
  wire multm_reduce_mulb1_cq141;
  wire multm_reduce_mulb1_cq142;
  wire multm_reduce_mulb1_cq143;
  wire multm_reduce_mulb1_cq144;
  wire multm_reduce_mulb1_cq145;
  wire multm_reduce_mulb1_cq146;
  wire multm_reduce_mulb1_cq147;
  wire multm_reduce_mulb1_cq148;
  wire multm_reduce_mulb1_cq149;
  wire multm_reduce_mulb1_cq150;
  wire multm_reduce_mulb1_cq151;
  wire multm_reduce_mulb1_cq152;
  wire multm_reduce_mulb1_cq153;
  wire multm_reduce_mulb1_cq154;
  wire multm_reduce_mulb1_cq155;
  wire multm_reduce_mulb1_cq156;
  wire multm_reduce_mulb1_cq157;
  wire multm_reduce_mulb1_cq158;
  wire multm_reduce_mulb1_cq159;
  wire multm_reduce_mulb1_cq160;
  wire multm_reduce_mulb1_cq161;
  wire multm_reduce_mulb1_cq162;
  wire multm_reduce_mulb1_cq163;
  wire multm_reduce_mulb1_cq164;
  wire multm_reduce_mulb1_cq165;
  wire multm_reduce_mulb1_cq166;
  wire multm_reduce_mulb1_cq167;
  wire multm_reduce_mulb1_cq168;
  wire multm_reduce_mulb1_cq169;
  wire multm_reduce_mulb1_cq170;
  wire multm_reduce_mulb1_cq171;
  wire multm_reduce_mulb1_cq172;
  wire multm_reduce_mulb1_cq173;
  wire multm_reduce_mulb1_cq174;
  wire multm_reduce_mulb1_cq175;
  wire multm_reduce_mulb1_cq176;
  wire multm_reduce_mulb1_cq177;
  wire multm_reduce_mulb1_cq178;
  wire multm_reduce_mulb1_cq179;
  wire multm_reduce_mulb1_cq180;
  wire multm_reduce_mulb1_cq181;
  wire multm_reduce_mulb1_cq182;
  wire multm_reduce_mulb1_pc0;
  wire multm_reduce_mulb1_pc1;
  wire multm_reduce_mulb1_pc2;
  wire multm_reduce_mulb1_pc3;
  wire multm_reduce_mulb1_pc4;
  wire multm_reduce_mulb1_pc5;
  wire multm_reduce_mulb1_pc6;
  wire multm_reduce_mulb1_pc7;
  wire multm_reduce_mulb1_pc8;
  wire multm_reduce_mulb1_pc9;
  wire multm_reduce_mulb1_pc10;
  wire multm_reduce_mulb1_pc11;
  wire multm_reduce_mulb1_pc12;
  wire multm_reduce_mulb1_pc13;
  wire multm_reduce_mulb1_pc14;
  wire multm_reduce_mulb1_pc15;
  wire multm_reduce_mulb1_pc16;
  wire multm_reduce_mulb1_pc17;
  wire multm_reduce_mulb1_pc18;
  wire multm_reduce_mulb1_pc19;
  wire multm_reduce_mulb1_pc20;
  wire multm_reduce_mulb1_pc21;
  wire multm_reduce_mulb1_pc22;
  wire multm_reduce_mulb1_pc23;
  wire multm_reduce_mulb1_pc24;
  wire multm_reduce_mulb1_pc25;
  wire multm_reduce_mulb1_pc26;
  wire multm_reduce_mulb1_pc27;
  wire multm_reduce_mulb1_pc28;
  wire multm_reduce_mulb1_pc29;
  wire multm_reduce_mulb1_pc30;
  wire multm_reduce_mulb1_pc31;
  wire multm_reduce_mulb1_pc32;
  wire multm_reduce_mulb1_pc33;
  wire multm_reduce_mulb1_pc34;
  wire multm_reduce_mulb1_pc35;
  wire multm_reduce_mulb1_pc36;
  wire multm_reduce_mulb1_pc37;
  wire multm_reduce_mulb1_pc38;
  wire multm_reduce_mulb1_pc39;
  wire multm_reduce_mulb1_pc40;
  wire multm_reduce_mulb1_pc41;
  wire multm_reduce_mulb1_pc42;
  wire multm_reduce_mulb1_pc43;
  wire multm_reduce_mulb1_pc44;
  wire multm_reduce_mulb1_pc45;
  wire multm_reduce_mulb1_pc46;
  wire multm_reduce_mulb1_pc47;
  wire multm_reduce_mulb1_pc48;
  wire multm_reduce_mulb1_pc49;
  wire multm_reduce_mulb1_pc50;
  wire multm_reduce_mulb1_pc51;
  wire multm_reduce_mulb1_pc52;
  wire multm_reduce_mulb1_pc53;
  wire multm_reduce_mulb1_pc54;
  wire multm_reduce_mulb1_pc55;
  wire multm_reduce_mulb1_pc56;
  wire multm_reduce_mulb1_pc57;
  wire multm_reduce_mulb1_pc58;
  wire multm_reduce_mulb1_pc59;
  wire multm_reduce_mulb1_pc60;
  wire multm_reduce_mulb1_pc61;
  wire multm_reduce_mulb1_pc62;
  wire multm_reduce_mulb1_pc63;
  wire multm_reduce_mulb1_pc64;
  wire multm_reduce_mulb1_pc65;
  wire multm_reduce_mulb1_pc66;
  wire multm_reduce_mulb1_pc67;
  wire multm_reduce_mulb1_pc68;
  wire multm_reduce_mulb1_pc69;
  wire multm_reduce_mulb1_pc70;
  wire multm_reduce_mulb1_pc71;
  wire multm_reduce_mulb1_pc72;
  wire multm_reduce_mulb1_pc73;
  wire multm_reduce_mulb1_pc74;
  wire multm_reduce_mulb1_pc75;
  wire multm_reduce_mulb1_pc76;
  wire multm_reduce_mulb1_pc77;
  wire multm_reduce_mulb1_pc78;
  wire multm_reduce_mulb1_pc79;
  wire multm_reduce_mulb1_pc80;
  wire multm_reduce_mulb1_pc81;
  wire multm_reduce_mulb1_pc82;
  wire multm_reduce_mulb1_pc83;
  wire multm_reduce_mulb1_pc84;
  wire multm_reduce_mulb1_pc85;
  wire multm_reduce_mulb1_pc86;
  wire multm_reduce_mulb1_pc87;
  wire multm_reduce_mulb1_pc88;
  wire multm_reduce_mulb1_pc89;
  wire multm_reduce_mulb1_pc90;
  wire multm_reduce_mulb1_pc91;
  wire multm_reduce_mulb1_pc92;
  wire multm_reduce_mulb1_pc93;
  wire multm_reduce_mulb1_pc94;
  wire multm_reduce_mulb1_pc95;
  wire multm_reduce_mulb1_pc96;
  wire multm_reduce_mulb1_pc97;
  wire multm_reduce_mulb1_pc98;
  wire multm_reduce_mulb1_pc99;
  wire multm_reduce_mulb1_pc100;
  wire multm_reduce_mulb1_pc101;
  wire multm_reduce_mulb1_pc102;
  wire multm_reduce_mulb1_pc103;
  wire multm_reduce_mulb1_pc104;
  wire multm_reduce_mulb1_pc105;
  wire multm_reduce_mulb1_pc106;
  wire multm_reduce_mulb1_pc107;
  wire multm_reduce_mulb1_pc108;
  wire multm_reduce_mulb1_pc109;
  wire multm_reduce_mulb1_pc110;
  wire multm_reduce_mulb1_pc111;
  wire multm_reduce_mulb1_pc112;
  wire multm_reduce_mulb1_pc113;
  wire multm_reduce_mulb1_pc114;
  wire multm_reduce_mulb1_pc115;
  wire multm_reduce_mulb1_pc116;
  wire multm_reduce_mulb1_pc117;
  wire multm_reduce_mulb1_pc118;
  wire multm_reduce_mulb1_pc119;
  wire multm_reduce_mulb1_pc120;
  wire multm_reduce_mulb1_pc121;
  wire multm_reduce_mulb1_pc122;
  wire multm_reduce_mulb1_pc123;
  wire multm_reduce_mulb1_pc124;
  wire multm_reduce_mulb1_pc125;
  wire multm_reduce_mulb1_pc126;
  wire multm_reduce_mulb1_pc127;
  wire multm_reduce_mulb1_pc128;
  wire multm_reduce_mulb1_pc129;
  wire multm_reduce_mulb1_pc130;
  wire multm_reduce_mulb1_pc131;
  wire multm_reduce_mulb1_pc132;
  wire multm_reduce_mulb1_pc133;
  wire multm_reduce_mulb1_pc134;
  wire multm_reduce_mulb1_pc135;
  wire multm_reduce_mulb1_pc136;
  wire multm_reduce_mulb1_pc137;
  wire multm_reduce_mulb1_pc138;
  wire multm_reduce_mulb1_pc139;
  wire multm_reduce_mulb1_pc140;
  wire multm_reduce_mulb1_pc141;
  wire multm_reduce_mulb1_pc142;
  wire multm_reduce_mulb1_pc143;
  wire multm_reduce_mulb1_pc144;
  wire multm_reduce_mulb1_pc145;
  wire multm_reduce_mulb1_pc146;
  wire multm_reduce_mulb1_pc147;
  wire multm_reduce_mulb1_pc148;
  wire multm_reduce_mulb1_pc149;
  wire multm_reduce_mulb1_pc150;
  wire multm_reduce_mulb1_pc151;
  wire multm_reduce_mulb1_pc152;
  wire multm_reduce_mulb1_pc153;
  wire multm_reduce_mulb1_pc154;
  wire multm_reduce_mulb1_pc155;
  wire multm_reduce_mulb1_pc156;
  wire multm_reduce_mulb1_pc157;
  wire multm_reduce_mulb1_pc158;
  wire multm_reduce_mulb1_pc159;
  wire multm_reduce_mulb1_pc160;
  wire multm_reduce_mulb1_pc161;
  wire multm_reduce_mulb1_pc162;
  wire multm_reduce_mulb1_pc163;
  wire multm_reduce_mulb1_pc164;
  wire multm_reduce_mulb1_pc165;
  wire multm_reduce_mulb1_pc166;
  wire multm_reduce_mulb1_pc167;
  wire multm_reduce_mulb1_pc168;
  wire multm_reduce_mulb1_pc169;
  wire multm_reduce_mulb1_pc170;
  wire multm_reduce_mulb1_pc171;
  wire multm_reduce_mulb1_pc172;
  wire multm_reduce_mulb1_pc173;
  wire multm_reduce_mulb1_pc174;
  wire multm_reduce_mulb1_pc175;
  wire multm_reduce_mulb1_pc176;
  wire multm_reduce_mulb1_pc177;
  wire multm_reduce_mulb1_pc178;
  wire multm_reduce_mulb1_pc179;
  wire multm_reduce_mulb1_pc180;
  wire multm_reduce_mulb1_pc181;
  wire multm_reduce_mulb1_pc182;
  wire multm_reduce_mulb1_ps0;
  wire multm_reduce_mulb1_ps1;
  wire multm_reduce_mulb1_ps2;
  wire multm_reduce_mulb1_ps3;
  wire multm_reduce_mulb1_ps4;
  wire multm_reduce_mulb1_ps5;
  wire multm_reduce_mulb1_ps6;
  wire multm_reduce_mulb1_ps7;
  wire multm_reduce_mulb1_ps8;
  wire multm_reduce_mulb1_ps9;
  wire multm_reduce_mulb1_ps10;
  wire multm_reduce_mulb1_ps11;
  wire multm_reduce_mulb1_ps12;
  wire multm_reduce_mulb1_ps13;
  wire multm_reduce_mulb1_ps14;
  wire multm_reduce_mulb1_ps15;
  wire multm_reduce_mulb1_ps16;
  wire multm_reduce_mulb1_ps17;
  wire multm_reduce_mulb1_ps18;
  wire multm_reduce_mulb1_ps19;
  wire multm_reduce_mulb1_ps20;
  wire multm_reduce_mulb1_ps21;
  wire multm_reduce_mulb1_ps22;
  wire multm_reduce_mulb1_ps23;
  wire multm_reduce_mulb1_ps24;
  wire multm_reduce_mulb1_ps25;
  wire multm_reduce_mulb1_ps26;
  wire multm_reduce_mulb1_ps27;
  wire multm_reduce_mulb1_ps28;
  wire multm_reduce_mulb1_ps29;
  wire multm_reduce_mulb1_ps30;
  wire multm_reduce_mulb1_ps31;
  wire multm_reduce_mulb1_ps32;
  wire multm_reduce_mulb1_ps33;
  wire multm_reduce_mulb1_ps34;
  wire multm_reduce_mulb1_ps35;
  wire multm_reduce_mulb1_ps36;
  wire multm_reduce_mulb1_ps37;
  wire multm_reduce_mulb1_ps38;
  wire multm_reduce_mulb1_ps39;
  wire multm_reduce_mulb1_ps40;
  wire multm_reduce_mulb1_ps41;
  wire multm_reduce_mulb1_ps42;
  wire multm_reduce_mulb1_ps43;
  wire multm_reduce_mulb1_ps44;
  wire multm_reduce_mulb1_ps45;
  wire multm_reduce_mulb1_ps46;
  wire multm_reduce_mulb1_ps47;
  wire multm_reduce_mulb1_ps48;
  wire multm_reduce_mulb1_ps49;
  wire multm_reduce_mulb1_ps50;
  wire multm_reduce_mulb1_ps51;
  wire multm_reduce_mulb1_ps52;
  wire multm_reduce_mulb1_ps53;
  wire multm_reduce_mulb1_ps54;
  wire multm_reduce_mulb1_ps55;
  wire multm_reduce_mulb1_ps56;
  wire multm_reduce_mulb1_ps57;
  wire multm_reduce_mulb1_ps58;
  wire multm_reduce_mulb1_ps59;
  wire multm_reduce_mulb1_ps60;
  wire multm_reduce_mulb1_ps61;
  wire multm_reduce_mulb1_ps62;
  wire multm_reduce_mulb1_ps63;
  wire multm_reduce_mulb1_ps64;
  wire multm_reduce_mulb1_ps65;
  wire multm_reduce_mulb1_ps66;
  wire multm_reduce_mulb1_ps67;
  wire multm_reduce_mulb1_ps68;
  wire multm_reduce_mulb1_ps69;
  wire multm_reduce_mulb1_ps70;
  wire multm_reduce_mulb1_ps71;
  wire multm_reduce_mulb1_ps72;
  wire multm_reduce_mulb1_ps73;
  wire multm_reduce_mulb1_ps74;
  wire multm_reduce_mulb1_ps75;
  wire multm_reduce_mulb1_ps76;
  wire multm_reduce_mulb1_ps77;
  wire multm_reduce_mulb1_ps78;
  wire multm_reduce_mulb1_ps79;
  wire multm_reduce_mulb1_ps80;
  wire multm_reduce_mulb1_ps81;
  wire multm_reduce_mulb1_ps82;
  wire multm_reduce_mulb1_ps83;
  wire multm_reduce_mulb1_ps84;
  wire multm_reduce_mulb1_ps85;
  wire multm_reduce_mulb1_ps86;
  wire multm_reduce_mulb1_ps87;
  wire multm_reduce_mulb1_ps88;
  wire multm_reduce_mulb1_ps89;
  wire multm_reduce_mulb1_ps90;
  wire multm_reduce_mulb1_ps91;
  wire multm_reduce_mulb1_ps92;
  wire multm_reduce_mulb1_ps93;
  wire multm_reduce_mulb1_ps94;
  wire multm_reduce_mulb1_ps95;
  wire multm_reduce_mulb1_ps96;
  wire multm_reduce_mulb1_ps97;
  wire multm_reduce_mulb1_ps98;
  wire multm_reduce_mulb1_ps99;
  wire multm_reduce_mulb1_ps100;
  wire multm_reduce_mulb1_ps101;
  wire multm_reduce_mulb1_ps102;
  wire multm_reduce_mulb1_ps103;
  wire multm_reduce_mulb1_ps104;
  wire multm_reduce_mulb1_ps105;
  wire multm_reduce_mulb1_ps106;
  wire multm_reduce_mulb1_ps107;
  wire multm_reduce_mulb1_ps108;
  wire multm_reduce_mulb1_ps109;
  wire multm_reduce_mulb1_ps110;
  wire multm_reduce_mulb1_ps111;
  wire multm_reduce_mulb1_ps112;
  wire multm_reduce_mulb1_ps113;
  wire multm_reduce_mulb1_ps114;
  wire multm_reduce_mulb1_ps115;
  wire multm_reduce_mulb1_ps116;
  wire multm_reduce_mulb1_ps117;
  wire multm_reduce_mulb1_ps118;
  wire multm_reduce_mulb1_ps119;
  wire multm_reduce_mulb1_ps120;
  wire multm_reduce_mulb1_ps121;
  wire multm_reduce_mulb1_ps122;
  wire multm_reduce_mulb1_ps123;
  wire multm_reduce_mulb1_ps124;
  wire multm_reduce_mulb1_ps125;
  wire multm_reduce_mulb1_ps126;
  wire multm_reduce_mulb1_ps127;
  wire multm_reduce_mulb1_ps128;
  wire multm_reduce_mulb1_ps129;
  wire multm_reduce_mulb1_ps130;
  wire multm_reduce_mulb1_ps131;
  wire multm_reduce_mulb1_ps132;
  wire multm_reduce_mulb1_ps133;
  wire multm_reduce_mulb1_ps134;
  wire multm_reduce_mulb1_ps135;
  wire multm_reduce_mulb1_ps136;
  wire multm_reduce_mulb1_ps137;
  wire multm_reduce_mulb1_ps138;
  wire multm_reduce_mulb1_ps139;
  wire multm_reduce_mulb1_ps140;
  wire multm_reduce_mulb1_ps141;
  wire multm_reduce_mulb1_ps142;
  wire multm_reduce_mulb1_ps143;
  wire multm_reduce_mulb1_ps144;
  wire multm_reduce_mulb1_ps145;
  wire multm_reduce_mulb1_ps146;
  wire multm_reduce_mulb1_ps147;
  wire multm_reduce_mulb1_ps148;
  wire multm_reduce_mulb1_ps149;
  wire multm_reduce_mulb1_ps150;
  wire multm_reduce_mulb1_ps151;
  wire multm_reduce_mulb1_ps152;
  wire multm_reduce_mulb1_ps153;
  wire multm_reduce_mulb1_ps154;
  wire multm_reduce_mulb1_ps155;
  wire multm_reduce_mulb1_ps156;
  wire multm_reduce_mulb1_ps157;
  wire multm_reduce_mulb1_ps158;
  wire multm_reduce_mulb1_ps159;
  wire multm_reduce_mulb1_ps160;
  wire multm_reduce_mulb1_ps161;
  wire multm_reduce_mulb1_ps162;
  wire multm_reduce_mulb1_ps163;
  wire multm_reduce_mulb1_ps164;
  wire multm_reduce_mulb1_ps165;
  wire multm_reduce_mulb1_ps166;
  wire multm_reduce_mulb1_ps167;
  wire multm_reduce_mulb1_ps168;
  wire multm_reduce_mulb1_ps169;
  wire multm_reduce_mulb1_ps170;
  wire multm_reduce_mulb1_ps171;
  wire multm_reduce_mulb1_ps172;
  wire multm_reduce_mulb1_ps173;
  wire multm_reduce_mulb1_ps174;
  wire multm_reduce_mulb1_ps175;
  wire multm_reduce_mulb1_ps176;
  wire multm_reduce_mulb1_ps177;
  wire multm_reduce_mulb1_ps178;
  wire multm_reduce_mulb1_ps179;
  wire multm_reduce_mulb1_ps180;
  wire multm_reduce_mulb1_ps181;
  wire multm_reduce_mulb1_sq0;
  wire multm_reduce_mulb1_sq1;
  wire multm_reduce_mulb1_sq2;
  wire multm_reduce_mulb1_sq3;
  wire multm_reduce_mulb1_sq4;
  wire multm_reduce_mulb1_sq5;
  wire multm_reduce_mulb1_sq6;
  wire multm_reduce_mulb1_sq7;
  wire multm_reduce_mulb1_sq8;
  wire multm_reduce_mulb1_sq9;
  wire multm_reduce_mulb1_sq10;
  wire multm_reduce_mulb1_sq11;
  wire multm_reduce_mulb1_sq12;
  wire multm_reduce_mulb1_sq13;
  wire multm_reduce_mulb1_sq14;
  wire multm_reduce_mulb1_sq15;
  wire multm_reduce_mulb1_sq16;
  wire multm_reduce_mulb1_sq17;
  wire multm_reduce_mulb1_sq18;
  wire multm_reduce_mulb1_sq19;
  wire multm_reduce_mulb1_sq20;
  wire multm_reduce_mulb1_sq21;
  wire multm_reduce_mulb1_sq22;
  wire multm_reduce_mulb1_sq23;
  wire multm_reduce_mulb1_sq24;
  wire multm_reduce_mulb1_sq25;
  wire multm_reduce_mulb1_sq26;
  wire multm_reduce_mulb1_sq27;
  wire multm_reduce_mulb1_sq28;
  wire multm_reduce_mulb1_sq29;
  wire multm_reduce_mulb1_sq30;
  wire multm_reduce_mulb1_sq31;
  wire multm_reduce_mulb1_sq32;
  wire multm_reduce_mulb1_sq33;
  wire multm_reduce_mulb1_sq34;
  wire multm_reduce_mulb1_sq35;
  wire multm_reduce_mulb1_sq36;
  wire multm_reduce_mulb1_sq37;
  wire multm_reduce_mulb1_sq38;
  wire multm_reduce_mulb1_sq39;
  wire multm_reduce_mulb1_sq40;
  wire multm_reduce_mulb1_sq41;
  wire multm_reduce_mulb1_sq42;
  wire multm_reduce_mulb1_sq43;
  wire multm_reduce_mulb1_sq44;
  wire multm_reduce_mulb1_sq45;
  wire multm_reduce_mulb1_sq46;
  wire multm_reduce_mulb1_sq47;
  wire multm_reduce_mulb1_sq48;
  wire multm_reduce_mulb1_sq49;
  wire multm_reduce_mulb1_sq50;
  wire multm_reduce_mulb1_sq51;
  wire multm_reduce_mulb1_sq52;
  wire multm_reduce_mulb1_sq53;
  wire multm_reduce_mulb1_sq54;
  wire multm_reduce_mulb1_sq55;
  wire multm_reduce_mulb1_sq56;
  wire multm_reduce_mulb1_sq57;
  wire multm_reduce_mulb1_sq58;
  wire multm_reduce_mulb1_sq59;
  wire multm_reduce_mulb1_sq60;
  wire multm_reduce_mulb1_sq61;
  wire multm_reduce_mulb1_sq62;
  wire multm_reduce_mulb1_sq63;
  wire multm_reduce_mulb1_sq64;
  wire multm_reduce_mulb1_sq65;
  wire multm_reduce_mulb1_sq66;
  wire multm_reduce_mulb1_sq67;
  wire multm_reduce_mulb1_sq68;
  wire multm_reduce_mulb1_sq69;
  wire multm_reduce_mulb1_sq70;
  wire multm_reduce_mulb1_sq71;
  wire multm_reduce_mulb1_sq72;
  wire multm_reduce_mulb1_sq73;
  wire multm_reduce_mulb1_sq74;
  wire multm_reduce_mulb1_sq75;
  wire multm_reduce_mulb1_sq76;
  wire multm_reduce_mulb1_sq77;
  wire multm_reduce_mulb1_sq78;
  wire multm_reduce_mulb1_sq79;
  wire multm_reduce_mulb1_sq80;
  wire multm_reduce_mulb1_sq81;
  wire multm_reduce_mulb1_sq82;
  wire multm_reduce_mulb1_sq83;
  wire multm_reduce_mulb1_sq84;
  wire multm_reduce_mulb1_sq85;
  wire multm_reduce_mulb1_sq86;
  wire multm_reduce_mulb1_sq87;
  wire multm_reduce_mulb1_sq88;
  wire multm_reduce_mulb1_sq89;
  wire multm_reduce_mulb1_sq90;
  wire multm_reduce_mulb1_sq91;
  wire multm_reduce_mulb1_sq92;
  wire multm_reduce_mulb1_sq93;
  wire multm_reduce_mulb1_sq94;
  wire multm_reduce_mulb1_sq95;
  wire multm_reduce_mulb1_sq96;
  wire multm_reduce_mulb1_sq97;
  wire multm_reduce_mulb1_sq98;
  wire multm_reduce_mulb1_sq99;
  wire multm_reduce_mulb1_sq100;
  wire multm_reduce_mulb1_sq101;
  wire multm_reduce_mulb1_sq102;
  wire multm_reduce_mulb1_sq103;
  wire multm_reduce_mulb1_sq104;
  wire multm_reduce_mulb1_sq105;
  wire multm_reduce_mulb1_sq106;
  wire multm_reduce_mulb1_sq107;
  wire multm_reduce_mulb1_sq108;
  wire multm_reduce_mulb1_sq109;
  wire multm_reduce_mulb1_sq110;
  wire multm_reduce_mulb1_sq111;
  wire multm_reduce_mulb1_sq112;
  wire multm_reduce_mulb1_sq113;
  wire multm_reduce_mulb1_sq114;
  wire multm_reduce_mulb1_sq115;
  wire multm_reduce_mulb1_sq116;
  wire multm_reduce_mulb1_sq117;
  wire multm_reduce_mulb1_sq118;
  wire multm_reduce_mulb1_sq119;
  wire multm_reduce_mulb1_sq120;
  wire multm_reduce_mulb1_sq121;
  wire multm_reduce_mulb1_sq122;
  wire multm_reduce_mulb1_sq123;
  wire multm_reduce_mulb1_sq124;
  wire multm_reduce_mulb1_sq125;
  wire multm_reduce_mulb1_sq126;
  wire multm_reduce_mulb1_sq127;
  wire multm_reduce_mulb1_sq128;
  wire multm_reduce_mulb1_sq129;
  wire multm_reduce_mulb1_sq130;
  wire multm_reduce_mulb1_sq131;
  wire multm_reduce_mulb1_sq132;
  wire multm_reduce_mulb1_sq133;
  wire multm_reduce_mulb1_sq134;
  wire multm_reduce_mulb1_sq135;
  wire multm_reduce_mulb1_sq136;
  wire multm_reduce_mulb1_sq137;
  wire multm_reduce_mulb1_sq138;
  wire multm_reduce_mulb1_sq139;
  wire multm_reduce_mulb1_sq140;
  wire multm_reduce_mulb1_sq141;
  wire multm_reduce_mulb1_sq142;
  wire multm_reduce_mulb1_sq143;
  wire multm_reduce_mulb1_sq144;
  wire multm_reduce_mulb1_sq145;
  wire multm_reduce_mulb1_sq146;
  wire multm_reduce_mulb1_sq147;
  wire multm_reduce_mulb1_sq148;
  wire multm_reduce_mulb1_sq149;
  wire multm_reduce_mulb1_sq150;
  wire multm_reduce_mulb1_sq151;
  wire multm_reduce_mulb1_sq152;
  wire multm_reduce_mulb1_sq153;
  wire multm_reduce_mulb1_sq154;
  wire multm_reduce_mulb1_sq155;
  wire multm_reduce_mulb1_sq156;
  wire multm_reduce_mulb1_sq157;
  wire multm_reduce_mulb1_sq158;
  wire multm_reduce_mulb1_sq159;
  wire multm_reduce_mulb1_sq160;
  wire multm_reduce_mulb1_sq161;
  wire multm_reduce_mulb1_sq162;
  wire multm_reduce_mulb1_sq163;
  wire multm_reduce_mulb1_sq164;
  wire multm_reduce_mulb1_sq165;
  wire multm_reduce_mulb1_sq166;
  wire multm_reduce_mulb1_sq167;
  wire multm_reduce_mulb1_sq168;
  wire multm_reduce_mulb1_sq169;
  wire multm_reduce_mulb1_sq170;
  wire multm_reduce_mulb1_sq171;
  wire multm_reduce_mulb1_sq172;
  wire multm_reduce_mulb1_sq173;
  wire multm_reduce_mulb1_sq174;
  wire multm_reduce_mulb1_sq175;
  wire multm_reduce_mulb1_sq176;
  wire multm_reduce_mulb1_sq177;
  wire multm_reduce_mulb1_sq178;
  wire multm_reduce_mulb1_sq179;
  wire multm_reduce_mulb1_sq180;
  wire multm_reduce_mulb1_sq181;
  wire multm_reduce_mulb1_sq182;
  wire multm_reduce_mulsc_mulb_add3_maj3_or3_wx;
  wire multm_reduce_mulsc_mulb_add3_maj3_wx;
  wire multm_reduce_mulsc_mulb_add3_maj3_wy;
  wire multm_reduce_mulsc_mulb_add3_maj3_xy;
  wire multm_reduce_mulsc_mulb_add3_xor3_wx;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx0;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx1;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx2;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx3;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx4;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx5;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx6;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx7;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx8;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx9;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx10;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx11;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx12;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx13;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx14;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx15;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx16;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx17;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx18;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx19;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx20;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx21;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx22;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx23;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx24;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx25;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx26;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx27;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx28;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx29;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx30;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx31;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx32;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx33;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx34;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx35;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx36;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx37;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx38;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx39;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx40;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx41;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx42;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx43;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx44;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx45;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx46;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx47;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx48;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx49;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx50;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx51;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx52;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx53;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx54;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx55;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx56;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx57;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx58;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx59;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx60;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx61;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx62;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx63;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx64;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx65;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx66;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx67;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx68;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx69;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx70;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx71;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx72;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx73;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx74;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx75;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx76;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx77;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx78;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx79;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx80;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx81;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx82;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx83;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx84;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx85;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx86;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx87;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx88;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx89;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx90;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx91;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx92;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx93;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx94;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx95;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx96;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx97;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx98;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx99;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx100;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx101;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx102;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx103;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx104;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx105;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx106;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx107;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx108;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx109;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx110;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx111;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx112;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx113;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx114;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx115;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx116;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx117;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx118;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx119;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx120;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx121;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx122;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx123;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx124;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx125;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx126;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx127;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx128;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx129;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx130;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx131;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx132;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx133;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx134;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx135;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx136;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx137;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx138;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx139;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx140;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx141;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx142;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx143;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx144;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx145;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx146;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx147;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx148;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx149;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx150;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx151;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx152;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx153;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx154;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx155;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx156;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx157;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx158;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx159;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx160;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx161;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx162;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx163;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx164;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx165;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx166;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx167;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx168;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx169;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx170;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx171;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx172;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx173;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx174;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx175;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx176;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx177;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx178;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx179;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx180;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx181;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx182;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx0;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx1;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx2;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx3;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx4;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx5;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx6;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx7;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx8;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx9;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx10;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx11;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx12;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx13;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx14;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx15;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx16;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx17;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx18;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx19;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx20;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx21;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx22;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx23;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx24;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx25;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx26;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx27;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx28;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx29;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx30;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx31;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx32;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx33;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx34;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx35;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx36;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx37;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx38;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx39;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx40;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx41;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx42;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx43;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx44;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx45;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx46;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx47;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx48;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx49;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx50;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx51;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx52;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx53;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx54;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx55;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx56;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx57;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx58;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx59;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx60;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx61;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx62;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx63;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx64;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx65;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx66;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx67;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx68;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx69;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx70;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx71;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx72;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx73;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx74;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx75;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx76;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx77;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx78;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx79;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx80;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx81;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx82;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx83;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx84;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx85;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx86;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx87;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx88;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx89;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx90;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx91;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx92;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx93;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx94;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx95;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx96;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx97;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx98;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx99;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx100;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx101;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx102;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx103;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx104;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx105;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx106;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx107;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx108;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx109;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx110;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx111;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx112;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx113;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx114;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx115;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx116;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx117;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx118;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx119;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx120;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx121;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx122;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx123;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx124;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx125;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx126;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx127;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx128;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx129;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx130;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx131;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx132;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx133;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx134;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx135;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx136;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx137;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx138;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx139;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx140;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx141;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx142;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx143;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx144;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx145;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx146;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx147;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx148;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx149;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx150;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx151;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx152;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx153;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx154;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx155;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx156;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx157;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx158;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx159;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx160;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx161;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx162;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx163;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx164;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx165;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx166;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx167;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx168;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx169;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx170;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx171;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx172;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx173;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx174;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx175;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx176;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx177;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx178;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx179;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx180;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx181;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wx182;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy0;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy1;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy2;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy3;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy4;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy5;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy6;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy7;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy8;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy9;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy10;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy11;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy12;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy13;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy14;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy15;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy16;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy17;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy18;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy19;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy20;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy21;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy22;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy23;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy24;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy25;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy26;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy27;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy28;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy29;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy30;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy31;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy32;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy33;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy34;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy35;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy36;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy37;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy38;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy39;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy40;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy41;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy42;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy43;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy44;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy45;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy46;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy47;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy48;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy49;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy50;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy51;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy52;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy53;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy54;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy55;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy56;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy57;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy58;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy59;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy60;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy61;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy62;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy63;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy64;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy65;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy66;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy67;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy68;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy69;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy70;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy71;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy72;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy73;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy74;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy75;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy76;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy77;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy78;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy79;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy80;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy81;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy82;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy83;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy84;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy85;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy86;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy87;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy88;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy89;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy90;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy91;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy92;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy93;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy94;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy95;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy96;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy97;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy98;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy99;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy100;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy101;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy102;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy103;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy104;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy105;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy106;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy107;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy108;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy109;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy110;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy111;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy112;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy113;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy114;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy115;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy116;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy117;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy118;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy119;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy120;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy121;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy122;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy123;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy124;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy125;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy126;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy127;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy128;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy129;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy130;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy131;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy132;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy133;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy134;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy135;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy136;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy137;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy138;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy139;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy140;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy141;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy142;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy143;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy144;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy145;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy146;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy147;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy148;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy149;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy150;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy151;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy152;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy153;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy154;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy155;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy156;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy157;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy158;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy159;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy160;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy161;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy162;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy163;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy164;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy165;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy166;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy167;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy168;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy169;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy170;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy171;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy172;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy173;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy174;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy175;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy176;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy177;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy178;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy179;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy180;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy181;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_wy182;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy0;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy1;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy2;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy3;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy4;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy5;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy6;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy7;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy8;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy9;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy10;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy11;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy12;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy13;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy14;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy15;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy16;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy17;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy18;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy19;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy20;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy21;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy22;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy23;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy24;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy25;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy26;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy27;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy28;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy29;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy30;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy31;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy32;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy33;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy34;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy35;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy36;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy37;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy38;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy39;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy40;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy41;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy42;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy43;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy44;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy45;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy46;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy47;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy48;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy49;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy50;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy51;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy52;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy53;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy54;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy55;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy56;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy57;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy58;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy59;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy60;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy61;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy62;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy63;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy64;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy65;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy66;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy67;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy68;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy69;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy70;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy71;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy72;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy73;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy74;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy75;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy76;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy77;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy78;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy79;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy80;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy81;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy82;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy83;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy84;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy85;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy86;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy87;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy88;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy89;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy90;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy91;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy92;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy93;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy94;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy95;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy96;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy97;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy98;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy99;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy100;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy101;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy102;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy103;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy104;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy105;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy106;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy107;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy108;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy109;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy110;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy111;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy112;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy113;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy114;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy115;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy116;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy117;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy118;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy119;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy120;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy121;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy122;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy123;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy124;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy125;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy126;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy127;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy128;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy129;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy130;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy131;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy132;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy133;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy134;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy135;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy136;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy137;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy138;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy139;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy140;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy141;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy142;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy143;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy144;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy145;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy146;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy147;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy148;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy149;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy150;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy151;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy152;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy153;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy154;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy155;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy156;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy157;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy158;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy159;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy160;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy161;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy162;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy163;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy164;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy165;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy166;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy167;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy168;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy169;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy170;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy171;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy172;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy173;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy174;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy175;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy176;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy177;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy178;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy179;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy180;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy181;
  wire multm_reduce_mulsc_mulb_add3b0_maj3b_xy182;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx0;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx1;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx2;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx3;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx4;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx5;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx6;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx7;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx8;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx9;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx10;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx11;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx12;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx13;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx14;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx15;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx16;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx17;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx18;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx19;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx20;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx21;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx22;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx23;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx24;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx25;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx26;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx27;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx28;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx29;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx30;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx31;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx32;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx33;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx34;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx35;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx36;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx37;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx38;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx39;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx40;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx41;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx42;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx43;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx44;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx45;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx46;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx47;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx48;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx49;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx50;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx51;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx52;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx53;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx54;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx55;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx56;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx57;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx58;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx59;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx60;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx61;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx62;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx63;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx64;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx65;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx66;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx67;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx68;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx69;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx70;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx71;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx72;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx73;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx74;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx75;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx76;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx77;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx78;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx79;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx80;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx81;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx82;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx83;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx84;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx85;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx86;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx87;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx88;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx89;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx90;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx91;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx92;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx93;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx94;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx95;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx96;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx97;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx98;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx99;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx100;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx101;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx102;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx103;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx104;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx105;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx106;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx107;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx108;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx109;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx110;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx111;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx112;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx113;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx114;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx115;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx116;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx117;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx118;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx119;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx120;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx121;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx122;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx123;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx124;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx125;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx126;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx127;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx128;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx129;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx130;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx131;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx132;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx133;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx134;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx135;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx136;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx137;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx138;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx139;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx140;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx141;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx142;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx143;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx144;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx145;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx146;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx147;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx148;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx149;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx150;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx151;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx152;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx153;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx154;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx155;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx156;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx157;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx158;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx159;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx160;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx161;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx162;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx163;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx164;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx165;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx166;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx167;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx168;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx169;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx170;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx171;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx172;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx173;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx174;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx175;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx176;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx177;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx178;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx179;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx180;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx181;
  wire multm_reduce_mulsc_mulb_add3b0_xor3b_wx182;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx0;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx1;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx2;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx3;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx4;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx5;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx6;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx7;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx8;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx9;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx10;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx11;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx12;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx13;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx14;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx15;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx16;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx17;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx18;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx19;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx20;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx21;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx22;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx23;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx24;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx25;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx26;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx27;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx28;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx29;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx30;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx31;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx32;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx33;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx34;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx35;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx36;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx37;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx38;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx39;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx40;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx41;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx42;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx43;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx44;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx45;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx46;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx47;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx48;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx49;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx50;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx51;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx52;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx53;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx54;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx55;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx56;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx57;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx58;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx59;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx60;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx61;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx62;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx63;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx64;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx65;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx66;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx67;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx68;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx69;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx70;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx71;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx72;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx73;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx74;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx75;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx76;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx77;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx78;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx79;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx80;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx81;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx82;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx83;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx84;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx85;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx86;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx87;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx88;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx89;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx90;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx91;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx92;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx93;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx94;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx95;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx96;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx97;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx98;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx99;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx100;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx101;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx102;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx103;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx104;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx105;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx106;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx107;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx108;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx109;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx110;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx111;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx112;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx113;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx114;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx115;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx116;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx117;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx118;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx119;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx120;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx121;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx122;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx123;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx124;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx125;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx126;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx127;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx128;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx129;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx130;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx131;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx132;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx133;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx134;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx135;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx136;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx137;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx138;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx139;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx140;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx141;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx142;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx143;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx144;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx145;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx146;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx147;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx148;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx149;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx150;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx151;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx152;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx153;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx154;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx155;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx156;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx157;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx158;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx159;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx160;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx161;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx162;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx163;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx164;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx165;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx166;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx167;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx168;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx169;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx170;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx171;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx172;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx173;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx174;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx175;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx176;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx177;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx178;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx179;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx180;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx181;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx182;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx0;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx1;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx2;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx3;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx4;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx5;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx6;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx7;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx8;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx9;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx10;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx11;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx12;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx13;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx14;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx15;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx16;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx17;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx18;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx19;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx20;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx21;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx22;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx23;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx24;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx25;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx26;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx27;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx28;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx29;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx30;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx31;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx32;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx33;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx34;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx35;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx36;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx37;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx38;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx39;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx40;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx41;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx42;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx43;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx44;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx45;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx46;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx47;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx48;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx49;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx50;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx51;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx52;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx53;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx54;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx55;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx56;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx57;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx58;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx59;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx60;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx61;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx62;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx63;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx64;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx65;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx66;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx67;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx68;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx69;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx70;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx71;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx72;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx73;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx74;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx75;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx76;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx77;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx78;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx79;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx80;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx81;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx82;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx83;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx84;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx85;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx86;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx87;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx88;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx89;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx90;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx91;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx92;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx93;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx94;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx95;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx96;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx97;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx98;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx99;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx100;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx101;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx102;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx103;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx104;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx105;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx106;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx107;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx108;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx109;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx110;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx111;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx112;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx113;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx114;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx115;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx116;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx117;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx118;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx119;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx120;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx121;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx122;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx123;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx124;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx125;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx126;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx127;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx128;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx129;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx130;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx131;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx132;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx133;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx134;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx135;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx136;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx137;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx138;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx139;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx140;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx141;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx142;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx143;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx144;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx145;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx146;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx147;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx148;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx149;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx150;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx151;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx152;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx153;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx154;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx155;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx156;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx157;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx158;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx159;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx160;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx161;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx162;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx163;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx164;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx165;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx166;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx167;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx168;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx169;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx170;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx171;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx172;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx173;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx174;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx175;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx176;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx177;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx178;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx179;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx180;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx181;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wx182;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy0;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy1;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy2;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy3;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy4;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy5;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy6;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy7;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy8;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy9;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy10;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy11;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy12;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy13;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy14;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy15;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy16;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy17;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy18;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy19;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy20;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy21;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy22;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy23;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy24;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy25;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy26;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy27;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy28;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy29;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy30;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy31;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy32;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy33;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy34;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy35;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy36;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy37;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy38;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy39;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy40;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy41;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy42;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy43;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy44;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy45;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy46;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy47;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy48;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy49;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy50;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy51;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy52;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy53;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy54;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy55;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy56;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy57;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy58;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy59;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy60;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy61;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy62;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy63;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy64;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy65;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy66;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy67;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy68;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy69;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy70;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy71;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy72;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy73;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy74;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy75;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy76;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy77;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy78;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy79;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy80;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy81;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy82;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy83;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy84;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy85;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy86;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy87;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy88;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy89;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy90;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy91;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy92;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy93;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy94;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy95;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy96;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy97;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy98;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy99;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy100;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy101;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy102;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy103;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy104;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy105;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy106;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy107;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy108;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy109;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy110;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy111;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy112;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy113;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy114;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy115;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy116;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy117;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy118;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy119;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy120;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy121;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy122;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy123;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy124;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy125;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy126;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy127;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy128;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy129;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy130;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy131;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy132;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy133;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy134;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy135;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy136;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy137;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy138;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy139;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy140;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy141;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy142;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy143;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy144;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy145;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy146;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy147;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy148;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy149;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy150;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy151;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy152;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy153;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy154;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy155;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy156;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy157;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy158;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy159;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy160;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy161;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy162;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy163;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy164;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy165;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy166;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy167;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy168;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy169;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy170;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy171;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy172;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy173;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy174;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy175;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy176;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy177;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy178;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy179;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy180;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy181;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_wy182;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy0;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy1;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy2;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy3;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy4;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy5;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy6;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy7;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy8;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy9;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy10;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy11;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy12;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy13;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy14;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy15;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy16;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy17;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy18;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy19;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy20;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy21;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy22;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy23;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy24;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy25;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy26;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy27;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy28;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy29;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy30;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy31;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy32;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy33;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy34;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy35;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy36;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy37;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy38;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy39;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy40;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy41;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy42;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy43;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy44;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy45;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy46;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy47;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy48;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy49;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy50;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy51;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy52;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy53;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy54;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy55;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy56;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy57;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy58;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy59;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy60;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy61;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy62;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy63;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy64;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy65;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy66;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy67;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy68;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy69;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy70;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy71;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy72;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy73;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy74;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy75;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy76;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy77;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy78;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy79;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy80;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy81;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy82;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy83;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy84;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy85;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy86;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy87;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy88;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy89;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy90;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy91;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy92;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy93;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy94;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy95;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy96;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy97;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy98;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy99;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy100;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy101;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy102;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy103;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy104;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy105;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy106;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy107;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy108;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy109;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy110;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy111;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy112;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy113;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy114;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy115;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy116;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy117;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy118;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy119;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy120;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy121;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy122;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy123;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy124;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy125;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy126;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy127;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy128;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy129;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy130;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy131;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy132;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy133;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy134;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy135;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy136;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy137;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy138;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy139;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy140;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy141;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy142;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy143;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy144;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy145;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy146;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy147;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy148;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy149;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy150;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy151;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy152;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy153;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy154;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy155;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy156;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy157;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy158;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy159;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy160;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy161;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy162;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy163;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy164;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy165;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy166;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy167;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy168;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy169;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy170;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy171;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy172;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy173;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy174;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy175;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy176;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy177;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy178;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy179;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy180;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy181;
  wire multm_reduce_mulsc_mulb_add3b1_maj3b_xy182;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx0;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx1;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx2;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx3;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx4;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx5;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx6;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx7;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx8;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx9;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx10;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx11;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx12;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx13;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx14;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx15;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx16;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx17;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx18;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx19;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx20;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx21;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx22;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx23;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx24;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx25;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx26;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx27;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx28;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx29;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx30;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx31;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx32;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx33;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx34;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx35;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx36;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx37;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx38;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx39;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx40;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx41;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx42;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx43;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx44;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx45;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx46;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx47;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx48;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx49;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx50;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx51;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx52;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx53;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx54;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx55;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx56;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx57;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx58;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx59;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx60;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx61;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx62;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx63;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx64;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx65;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx66;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx67;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx68;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx69;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx70;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx71;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx72;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx73;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx74;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx75;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx76;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx77;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx78;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx79;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx80;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx81;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx82;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx83;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx84;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx85;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx86;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx87;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx88;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx89;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx90;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx91;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx92;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx93;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx94;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx95;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx96;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx97;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx98;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx99;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx100;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx101;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx102;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx103;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx104;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx105;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx106;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx107;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx108;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx109;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx110;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx111;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx112;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx113;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx114;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx115;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx116;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx117;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx118;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx119;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx120;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx121;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx122;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx123;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx124;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx125;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx126;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx127;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx128;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx129;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx130;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx131;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx132;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx133;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx134;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx135;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx136;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx137;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx138;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx139;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx140;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx141;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx142;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx143;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx144;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx145;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx146;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx147;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx148;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx149;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx150;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx151;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx152;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx153;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx154;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx155;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx156;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx157;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx158;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx159;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx160;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx161;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx162;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx163;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx164;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx165;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx166;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx167;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx168;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx169;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx170;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx171;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx172;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx173;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx174;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx175;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx176;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx177;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx178;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx179;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx180;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx181;
  wire multm_reduce_mulsc_mulb_add3b1_xor3b_wx182;
  wire multm_reduce_mulsc_mulb_cq0;
  wire multm_reduce_mulsc_mulb_cq1;
  wire multm_reduce_mulsc_mulb_cq2;
  wire multm_reduce_mulsc_mulb_cq3;
  wire multm_reduce_mulsc_mulb_cq4;
  wire multm_reduce_mulsc_mulb_cq5;
  wire multm_reduce_mulsc_mulb_cq6;
  wire multm_reduce_mulsc_mulb_cq7;
  wire multm_reduce_mulsc_mulb_cq8;
  wire multm_reduce_mulsc_mulb_cq9;
  wire multm_reduce_mulsc_mulb_cq10;
  wire multm_reduce_mulsc_mulb_cq11;
  wire multm_reduce_mulsc_mulb_cq12;
  wire multm_reduce_mulsc_mulb_cq13;
  wire multm_reduce_mulsc_mulb_cq14;
  wire multm_reduce_mulsc_mulb_cq15;
  wire multm_reduce_mulsc_mulb_cq16;
  wire multm_reduce_mulsc_mulb_cq17;
  wire multm_reduce_mulsc_mulb_cq18;
  wire multm_reduce_mulsc_mulb_cq19;
  wire multm_reduce_mulsc_mulb_cq20;
  wire multm_reduce_mulsc_mulb_cq21;
  wire multm_reduce_mulsc_mulb_cq22;
  wire multm_reduce_mulsc_mulb_cq23;
  wire multm_reduce_mulsc_mulb_cq24;
  wire multm_reduce_mulsc_mulb_cq25;
  wire multm_reduce_mulsc_mulb_cq26;
  wire multm_reduce_mulsc_mulb_cq27;
  wire multm_reduce_mulsc_mulb_cq28;
  wire multm_reduce_mulsc_mulb_cq29;
  wire multm_reduce_mulsc_mulb_cq30;
  wire multm_reduce_mulsc_mulb_cq31;
  wire multm_reduce_mulsc_mulb_cq32;
  wire multm_reduce_mulsc_mulb_cq33;
  wire multm_reduce_mulsc_mulb_cq34;
  wire multm_reduce_mulsc_mulb_cq35;
  wire multm_reduce_mulsc_mulb_cq36;
  wire multm_reduce_mulsc_mulb_cq37;
  wire multm_reduce_mulsc_mulb_cq38;
  wire multm_reduce_mulsc_mulb_cq39;
  wire multm_reduce_mulsc_mulb_cq40;
  wire multm_reduce_mulsc_mulb_cq41;
  wire multm_reduce_mulsc_mulb_cq42;
  wire multm_reduce_mulsc_mulb_cq43;
  wire multm_reduce_mulsc_mulb_cq44;
  wire multm_reduce_mulsc_mulb_cq45;
  wire multm_reduce_mulsc_mulb_cq46;
  wire multm_reduce_mulsc_mulb_cq47;
  wire multm_reduce_mulsc_mulb_cq48;
  wire multm_reduce_mulsc_mulb_cq49;
  wire multm_reduce_mulsc_mulb_cq50;
  wire multm_reduce_mulsc_mulb_cq51;
  wire multm_reduce_mulsc_mulb_cq52;
  wire multm_reduce_mulsc_mulb_cq53;
  wire multm_reduce_mulsc_mulb_cq54;
  wire multm_reduce_mulsc_mulb_cq55;
  wire multm_reduce_mulsc_mulb_cq56;
  wire multm_reduce_mulsc_mulb_cq57;
  wire multm_reduce_mulsc_mulb_cq58;
  wire multm_reduce_mulsc_mulb_cq59;
  wire multm_reduce_mulsc_mulb_cq60;
  wire multm_reduce_mulsc_mulb_cq61;
  wire multm_reduce_mulsc_mulb_cq62;
  wire multm_reduce_mulsc_mulb_cq63;
  wire multm_reduce_mulsc_mulb_cq64;
  wire multm_reduce_mulsc_mulb_cq65;
  wire multm_reduce_mulsc_mulb_cq66;
  wire multm_reduce_mulsc_mulb_cq67;
  wire multm_reduce_mulsc_mulb_cq68;
  wire multm_reduce_mulsc_mulb_cq69;
  wire multm_reduce_mulsc_mulb_cq70;
  wire multm_reduce_mulsc_mulb_cq71;
  wire multm_reduce_mulsc_mulb_cq72;
  wire multm_reduce_mulsc_mulb_cq73;
  wire multm_reduce_mulsc_mulb_cq74;
  wire multm_reduce_mulsc_mulb_cq75;
  wire multm_reduce_mulsc_mulb_cq76;
  wire multm_reduce_mulsc_mulb_cq77;
  wire multm_reduce_mulsc_mulb_cq78;
  wire multm_reduce_mulsc_mulb_cq79;
  wire multm_reduce_mulsc_mulb_cq80;
  wire multm_reduce_mulsc_mulb_cq81;
  wire multm_reduce_mulsc_mulb_cq82;
  wire multm_reduce_mulsc_mulb_cq83;
  wire multm_reduce_mulsc_mulb_cq84;
  wire multm_reduce_mulsc_mulb_cq85;
  wire multm_reduce_mulsc_mulb_cq86;
  wire multm_reduce_mulsc_mulb_cq87;
  wire multm_reduce_mulsc_mulb_cq88;
  wire multm_reduce_mulsc_mulb_cq89;
  wire multm_reduce_mulsc_mulb_cq90;
  wire multm_reduce_mulsc_mulb_cq91;
  wire multm_reduce_mulsc_mulb_cq92;
  wire multm_reduce_mulsc_mulb_cq93;
  wire multm_reduce_mulsc_mulb_cq94;
  wire multm_reduce_mulsc_mulb_cq95;
  wire multm_reduce_mulsc_mulb_cq96;
  wire multm_reduce_mulsc_mulb_cq97;
  wire multm_reduce_mulsc_mulb_cq98;
  wire multm_reduce_mulsc_mulb_cq99;
  wire multm_reduce_mulsc_mulb_cq100;
  wire multm_reduce_mulsc_mulb_cq101;
  wire multm_reduce_mulsc_mulb_cq102;
  wire multm_reduce_mulsc_mulb_cq103;
  wire multm_reduce_mulsc_mulb_cq104;
  wire multm_reduce_mulsc_mulb_cq105;
  wire multm_reduce_mulsc_mulb_cq106;
  wire multm_reduce_mulsc_mulb_cq107;
  wire multm_reduce_mulsc_mulb_cq108;
  wire multm_reduce_mulsc_mulb_cq109;
  wire multm_reduce_mulsc_mulb_cq110;
  wire multm_reduce_mulsc_mulb_cq111;
  wire multm_reduce_mulsc_mulb_cq112;
  wire multm_reduce_mulsc_mulb_cq113;
  wire multm_reduce_mulsc_mulb_cq114;
  wire multm_reduce_mulsc_mulb_cq115;
  wire multm_reduce_mulsc_mulb_cq116;
  wire multm_reduce_mulsc_mulb_cq117;
  wire multm_reduce_mulsc_mulb_cq118;
  wire multm_reduce_mulsc_mulb_cq119;
  wire multm_reduce_mulsc_mulb_cq120;
  wire multm_reduce_mulsc_mulb_cq121;
  wire multm_reduce_mulsc_mulb_cq122;
  wire multm_reduce_mulsc_mulb_cq123;
  wire multm_reduce_mulsc_mulb_cq124;
  wire multm_reduce_mulsc_mulb_cq125;
  wire multm_reduce_mulsc_mulb_cq126;
  wire multm_reduce_mulsc_mulb_cq127;
  wire multm_reduce_mulsc_mulb_cq128;
  wire multm_reduce_mulsc_mulb_cq129;
  wire multm_reduce_mulsc_mulb_cq130;
  wire multm_reduce_mulsc_mulb_cq131;
  wire multm_reduce_mulsc_mulb_cq132;
  wire multm_reduce_mulsc_mulb_cq133;
  wire multm_reduce_mulsc_mulb_cq134;
  wire multm_reduce_mulsc_mulb_cq135;
  wire multm_reduce_mulsc_mulb_cq136;
  wire multm_reduce_mulsc_mulb_cq137;
  wire multm_reduce_mulsc_mulb_cq138;
  wire multm_reduce_mulsc_mulb_cq139;
  wire multm_reduce_mulsc_mulb_cq140;
  wire multm_reduce_mulsc_mulb_cq141;
  wire multm_reduce_mulsc_mulb_cq142;
  wire multm_reduce_mulsc_mulb_cq143;
  wire multm_reduce_mulsc_mulb_cq144;
  wire multm_reduce_mulsc_mulb_cq145;
  wire multm_reduce_mulsc_mulb_cq146;
  wire multm_reduce_mulsc_mulb_cq147;
  wire multm_reduce_mulsc_mulb_cq148;
  wire multm_reduce_mulsc_mulb_cq149;
  wire multm_reduce_mulsc_mulb_cq150;
  wire multm_reduce_mulsc_mulb_cq151;
  wire multm_reduce_mulsc_mulb_cq152;
  wire multm_reduce_mulsc_mulb_cq153;
  wire multm_reduce_mulsc_mulb_cq154;
  wire multm_reduce_mulsc_mulb_cq155;
  wire multm_reduce_mulsc_mulb_cq156;
  wire multm_reduce_mulsc_mulb_cq157;
  wire multm_reduce_mulsc_mulb_cq158;
  wire multm_reduce_mulsc_mulb_cq159;
  wire multm_reduce_mulsc_mulb_cq160;
  wire multm_reduce_mulsc_mulb_cq161;
  wire multm_reduce_mulsc_mulb_cq162;
  wire multm_reduce_mulsc_mulb_cq163;
  wire multm_reduce_mulsc_mulb_cq164;
  wire multm_reduce_mulsc_mulb_cq165;
  wire multm_reduce_mulsc_mulb_cq166;
  wire multm_reduce_mulsc_mulb_cq167;
  wire multm_reduce_mulsc_mulb_cq168;
  wire multm_reduce_mulsc_mulb_cq169;
  wire multm_reduce_mulsc_mulb_cq170;
  wire multm_reduce_mulsc_mulb_cq171;
  wire multm_reduce_mulsc_mulb_cq172;
  wire multm_reduce_mulsc_mulb_cq173;
  wire multm_reduce_mulsc_mulb_cq174;
  wire multm_reduce_mulsc_mulb_cq175;
  wire multm_reduce_mulsc_mulb_cq176;
  wire multm_reduce_mulsc_mulb_cq177;
  wire multm_reduce_mulsc_mulb_cq178;
  wire multm_reduce_mulsc_mulb_cq179;
  wire multm_reduce_mulsc_mulb_cq180;
  wire multm_reduce_mulsc_mulb_cq181;
  wire multm_reduce_mulsc_mulb_cq182;
  wire multm_reduce_mulsc_mulb_cq183;
  wire multm_reduce_mulsc_mulb_pc0;
  wire multm_reduce_mulsc_mulb_pc1;
  wire multm_reduce_mulsc_mulb_pc2;
  wire multm_reduce_mulsc_mulb_pc3;
  wire multm_reduce_mulsc_mulb_pc4;
  wire multm_reduce_mulsc_mulb_pc5;
  wire multm_reduce_mulsc_mulb_pc6;
  wire multm_reduce_mulsc_mulb_pc7;
  wire multm_reduce_mulsc_mulb_pc8;
  wire multm_reduce_mulsc_mulb_pc9;
  wire multm_reduce_mulsc_mulb_pc10;
  wire multm_reduce_mulsc_mulb_pc11;
  wire multm_reduce_mulsc_mulb_pc12;
  wire multm_reduce_mulsc_mulb_pc13;
  wire multm_reduce_mulsc_mulb_pc14;
  wire multm_reduce_mulsc_mulb_pc15;
  wire multm_reduce_mulsc_mulb_pc16;
  wire multm_reduce_mulsc_mulb_pc17;
  wire multm_reduce_mulsc_mulb_pc18;
  wire multm_reduce_mulsc_mulb_pc19;
  wire multm_reduce_mulsc_mulb_pc20;
  wire multm_reduce_mulsc_mulb_pc21;
  wire multm_reduce_mulsc_mulb_pc22;
  wire multm_reduce_mulsc_mulb_pc23;
  wire multm_reduce_mulsc_mulb_pc24;
  wire multm_reduce_mulsc_mulb_pc25;
  wire multm_reduce_mulsc_mulb_pc26;
  wire multm_reduce_mulsc_mulb_pc27;
  wire multm_reduce_mulsc_mulb_pc28;
  wire multm_reduce_mulsc_mulb_pc29;
  wire multm_reduce_mulsc_mulb_pc30;
  wire multm_reduce_mulsc_mulb_pc31;
  wire multm_reduce_mulsc_mulb_pc32;
  wire multm_reduce_mulsc_mulb_pc33;
  wire multm_reduce_mulsc_mulb_pc34;
  wire multm_reduce_mulsc_mulb_pc35;
  wire multm_reduce_mulsc_mulb_pc36;
  wire multm_reduce_mulsc_mulb_pc37;
  wire multm_reduce_mulsc_mulb_pc38;
  wire multm_reduce_mulsc_mulb_pc39;
  wire multm_reduce_mulsc_mulb_pc40;
  wire multm_reduce_mulsc_mulb_pc41;
  wire multm_reduce_mulsc_mulb_pc42;
  wire multm_reduce_mulsc_mulb_pc43;
  wire multm_reduce_mulsc_mulb_pc44;
  wire multm_reduce_mulsc_mulb_pc45;
  wire multm_reduce_mulsc_mulb_pc46;
  wire multm_reduce_mulsc_mulb_pc47;
  wire multm_reduce_mulsc_mulb_pc48;
  wire multm_reduce_mulsc_mulb_pc49;
  wire multm_reduce_mulsc_mulb_pc50;
  wire multm_reduce_mulsc_mulb_pc51;
  wire multm_reduce_mulsc_mulb_pc52;
  wire multm_reduce_mulsc_mulb_pc53;
  wire multm_reduce_mulsc_mulb_pc54;
  wire multm_reduce_mulsc_mulb_pc55;
  wire multm_reduce_mulsc_mulb_pc56;
  wire multm_reduce_mulsc_mulb_pc57;
  wire multm_reduce_mulsc_mulb_pc58;
  wire multm_reduce_mulsc_mulb_pc59;
  wire multm_reduce_mulsc_mulb_pc60;
  wire multm_reduce_mulsc_mulb_pc61;
  wire multm_reduce_mulsc_mulb_pc62;
  wire multm_reduce_mulsc_mulb_pc63;
  wire multm_reduce_mulsc_mulb_pc64;
  wire multm_reduce_mulsc_mulb_pc65;
  wire multm_reduce_mulsc_mulb_pc66;
  wire multm_reduce_mulsc_mulb_pc67;
  wire multm_reduce_mulsc_mulb_pc68;
  wire multm_reduce_mulsc_mulb_pc69;
  wire multm_reduce_mulsc_mulb_pc70;
  wire multm_reduce_mulsc_mulb_pc71;
  wire multm_reduce_mulsc_mulb_pc72;
  wire multm_reduce_mulsc_mulb_pc73;
  wire multm_reduce_mulsc_mulb_pc74;
  wire multm_reduce_mulsc_mulb_pc75;
  wire multm_reduce_mulsc_mulb_pc76;
  wire multm_reduce_mulsc_mulb_pc77;
  wire multm_reduce_mulsc_mulb_pc78;
  wire multm_reduce_mulsc_mulb_pc79;
  wire multm_reduce_mulsc_mulb_pc80;
  wire multm_reduce_mulsc_mulb_pc81;
  wire multm_reduce_mulsc_mulb_pc82;
  wire multm_reduce_mulsc_mulb_pc83;
  wire multm_reduce_mulsc_mulb_pc84;
  wire multm_reduce_mulsc_mulb_pc85;
  wire multm_reduce_mulsc_mulb_pc86;
  wire multm_reduce_mulsc_mulb_pc87;
  wire multm_reduce_mulsc_mulb_pc88;
  wire multm_reduce_mulsc_mulb_pc89;
  wire multm_reduce_mulsc_mulb_pc90;
  wire multm_reduce_mulsc_mulb_pc91;
  wire multm_reduce_mulsc_mulb_pc92;
  wire multm_reduce_mulsc_mulb_pc93;
  wire multm_reduce_mulsc_mulb_pc94;
  wire multm_reduce_mulsc_mulb_pc95;
  wire multm_reduce_mulsc_mulb_pc96;
  wire multm_reduce_mulsc_mulb_pc97;
  wire multm_reduce_mulsc_mulb_pc98;
  wire multm_reduce_mulsc_mulb_pc99;
  wire multm_reduce_mulsc_mulb_pc100;
  wire multm_reduce_mulsc_mulb_pc101;
  wire multm_reduce_mulsc_mulb_pc102;
  wire multm_reduce_mulsc_mulb_pc103;
  wire multm_reduce_mulsc_mulb_pc104;
  wire multm_reduce_mulsc_mulb_pc105;
  wire multm_reduce_mulsc_mulb_pc106;
  wire multm_reduce_mulsc_mulb_pc107;
  wire multm_reduce_mulsc_mulb_pc108;
  wire multm_reduce_mulsc_mulb_pc109;
  wire multm_reduce_mulsc_mulb_pc110;
  wire multm_reduce_mulsc_mulb_pc111;
  wire multm_reduce_mulsc_mulb_pc112;
  wire multm_reduce_mulsc_mulb_pc113;
  wire multm_reduce_mulsc_mulb_pc114;
  wire multm_reduce_mulsc_mulb_pc115;
  wire multm_reduce_mulsc_mulb_pc116;
  wire multm_reduce_mulsc_mulb_pc117;
  wire multm_reduce_mulsc_mulb_pc118;
  wire multm_reduce_mulsc_mulb_pc119;
  wire multm_reduce_mulsc_mulb_pc120;
  wire multm_reduce_mulsc_mulb_pc121;
  wire multm_reduce_mulsc_mulb_pc122;
  wire multm_reduce_mulsc_mulb_pc123;
  wire multm_reduce_mulsc_mulb_pc124;
  wire multm_reduce_mulsc_mulb_pc125;
  wire multm_reduce_mulsc_mulb_pc126;
  wire multm_reduce_mulsc_mulb_pc127;
  wire multm_reduce_mulsc_mulb_pc128;
  wire multm_reduce_mulsc_mulb_pc129;
  wire multm_reduce_mulsc_mulb_pc130;
  wire multm_reduce_mulsc_mulb_pc131;
  wire multm_reduce_mulsc_mulb_pc132;
  wire multm_reduce_mulsc_mulb_pc133;
  wire multm_reduce_mulsc_mulb_pc134;
  wire multm_reduce_mulsc_mulb_pc135;
  wire multm_reduce_mulsc_mulb_pc136;
  wire multm_reduce_mulsc_mulb_pc137;
  wire multm_reduce_mulsc_mulb_pc138;
  wire multm_reduce_mulsc_mulb_pc139;
  wire multm_reduce_mulsc_mulb_pc140;
  wire multm_reduce_mulsc_mulb_pc141;
  wire multm_reduce_mulsc_mulb_pc142;
  wire multm_reduce_mulsc_mulb_pc143;
  wire multm_reduce_mulsc_mulb_pc144;
  wire multm_reduce_mulsc_mulb_pc145;
  wire multm_reduce_mulsc_mulb_pc146;
  wire multm_reduce_mulsc_mulb_pc147;
  wire multm_reduce_mulsc_mulb_pc148;
  wire multm_reduce_mulsc_mulb_pc149;
  wire multm_reduce_mulsc_mulb_pc150;
  wire multm_reduce_mulsc_mulb_pc151;
  wire multm_reduce_mulsc_mulb_pc152;
  wire multm_reduce_mulsc_mulb_pc153;
  wire multm_reduce_mulsc_mulb_pc154;
  wire multm_reduce_mulsc_mulb_pc155;
  wire multm_reduce_mulsc_mulb_pc156;
  wire multm_reduce_mulsc_mulb_pc157;
  wire multm_reduce_mulsc_mulb_pc158;
  wire multm_reduce_mulsc_mulb_pc159;
  wire multm_reduce_mulsc_mulb_pc160;
  wire multm_reduce_mulsc_mulb_pc161;
  wire multm_reduce_mulsc_mulb_pc162;
  wire multm_reduce_mulsc_mulb_pc163;
  wire multm_reduce_mulsc_mulb_pc164;
  wire multm_reduce_mulsc_mulb_pc165;
  wire multm_reduce_mulsc_mulb_pc166;
  wire multm_reduce_mulsc_mulb_pc167;
  wire multm_reduce_mulsc_mulb_pc168;
  wire multm_reduce_mulsc_mulb_pc169;
  wire multm_reduce_mulsc_mulb_pc170;
  wire multm_reduce_mulsc_mulb_pc171;
  wire multm_reduce_mulsc_mulb_pc172;
  wire multm_reduce_mulsc_mulb_pc173;
  wire multm_reduce_mulsc_mulb_pc174;
  wire multm_reduce_mulsc_mulb_pc175;
  wire multm_reduce_mulsc_mulb_pc176;
  wire multm_reduce_mulsc_mulb_pc177;
  wire multm_reduce_mulsc_mulb_pc178;
  wire multm_reduce_mulsc_mulb_pc179;
  wire multm_reduce_mulsc_mulb_pc180;
  wire multm_reduce_mulsc_mulb_pc181;
  wire multm_reduce_mulsc_mulb_pc182;
  wire multm_reduce_mulsc_mulb_pc183;
  wire multm_reduce_mulsc_mulb_ps0;
  wire multm_reduce_mulsc_mulb_ps1;
  wire multm_reduce_mulsc_mulb_ps2;
  wire multm_reduce_mulsc_mulb_ps3;
  wire multm_reduce_mulsc_mulb_ps4;
  wire multm_reduce_mulsc_mulb_ps5;
  wire multm_reduce_mulsc_mulb_ps6;
  wire multm_reduce_mulsc_mulb_ps7;
  wire multm_reduce_mulsc_mulb_ps8;
  wire multm_reduce_mulsc_mulb_ps9;
  wire multm_reduce_mulsc_mulb_ps10;
  wire multm_reduce_mulsc_mulb_ps11;
  wire multm_reduce_mulsc_mulb_ps12;
  wire multm_reduce_mulsc_mulb_ps13;
  wire multm_reduce_mulsc_mulb_ps14;
  wire multm_reduce_mulsc_mulb_ps15;
  wire multm_reduce_mulsc_mulb_ps16;
  wire multm_reduce_mulsc_mulb_ps17;
  wire multm_reduce_mulsc_mulb_ps18;
  wire multm_reduce_mulsc_mulb_ps19;
  wire multm_reduce_mulsc_mulb_ps20;
  wire multm_reduce_mulsc_mulb_ps21;
  wire multm_reduce_mulsc_mulb_ps22;
  wire multm_reduce_mulsc_mulb_ps23;
  wire multm_reduce_mulsc_mulb_ps24;
  wire multm_reduce_mulsc_mulb_ps25;
  wire multm_reduce_mulsc_mulb_ps26;
  wire multm_reduce_mulsc_mulb_ps27;
  wire multm_reduce_mulsc_mulb_ps28;
  wire multm_reduce_mulsc_mulb_ps29;
  wire multm_reduce_mulsc_mulb_ps30;
  wire multm_reduce_mulsc_mulb_ps31;
  wire multm_reduce_mulsc_mulb_ps32;
  wire multm_reduce_mulsc_mulb_ps33;
  wire multm_reduce_mulsc_mulb_ps34;
  wire multm_reduce_mulsc_mulb_ps35;
  wire multm_reduce_mulsc_mulb_ps36;
  wire multm_reduce_mulsc_mulb_ps37;
  wire multm_reduce_mulsc_mulb_ps38;
  wire multm_reduce_mulsc_mulb_ps39;
  wire multm_reduce_mulsc_mulb_ps40;
  wire multm_reduce_mulsc_mulb_ps41;
  wire multm_reduce_mulsc_mulb_ps42;
  wire multm_reduce_mulsc_mulb_ps43;
  wire multm_reduce_mulsc_mulb_ps44;
  wire multm_reduce_mulsc_mulb_ps45;
  wire multm_reduce_mulsc_mulb_ps46;
  wire multm_reduce_mulsc_mulb_ps47;
  wire multm_reduce_mulsc_mulb_ps48;
  wire multm_reduce_mulsc_mulb_ps49;
  wire multm_reduce_mulsc_mulb_ps50;
  wire multm_reduce_mulsc_mulb_ps51;
  wire multm_reduce_mulsc_mulb_ps52;
  wire multm_reduce_mulsc_mulb_ps53;
  wire multm_reduce_mulsc_mulb_ps54;
  wire multm_reduce_mulsc_mulb_ps55;
  wire multm_reduce_mulsc_mulb_ps56;
  wire multm_reduce_mulsc_mulb_ps57;
  wire multm_reduce_mulsc_mulb_ps58;
  wire multm_reduce_mulsc_mulb_ps59;
  wire multm_reduce_mulsc_mulb_ps60;
  wire multm_reduce_mulsc_mulb_ps61;
  wire multm_reduce_mulsc_mulb_ps62;
  wire multm_reduce_mulsc_mulb_ps63;
  wire multm_reduce_mulsc_mulb_ps64;
  wire multm_reduce_mulsc_mulb_ps65;
  wire multm_reduce_mulsc_mulb_ps66;
  wire multm_reduce_mulsc_mulb_ps67;
  wire multm_reduce_mulsc_mulb_ps68;
  wire multm_reduce_mulsc_mulb_ps69;
  wire multm_reduce_mulsc_mulb_ps70;
  wire multm_reduce_mulsc_mulb_ps71;
  wire multm_reduce_mulsc_mulb_ps72;
  wire multm_reduce_mulsc_mulb_ps73;
  wire multm_reduce_mulsc_mulb_ps74;
  wire multm_reduce_mulsc_mulb_ps75;
  wire multm_reduce_mulsc_mulb_ps76;
  wire multm_reduce_mulsc_mulb_ps77;
  wire multm_reduce_mulsc_mulb_ps78;
  wire multm_reduce_mulsc_mulb_ps79;
  wire multm_reduce_mulsc_mulb_ps80;
  wire multm_reduce_mulsc_mulb_ps81;
  wire multm_reduce_mulsc_mulb_ps82;
  wire multm_reduce_mulsc_mulb_ps83;
  wire multm_reduce_mulsc_mulb_ps84;
  wire multm_reduce_mulsc_mulb_ps85;
  wire multm_reduce_mulsc_mulb_ps86;
  wire multm_reduce_mulsc_mulb_ps87;
  wire multm_reduce_mulsc_mulb_ps88;
  wire multm_reduce_mulsc_mulb_ps89;
  wire multm_reduce_mulsc_mulb_ps90;
  wire multm_reduce_mulsc_mulb_ps91;
  wire multm_reduce_mulsc_mulb_ps92;
  wire multm_reduce_mulsc_mulb_ps93;
  wire multm_reduce_mulsc_mulb_ps94;
  wire multm_reduce_mulsc_mulb_ps95;
  wire multm_reduce_mulsc_mulb_ps96;
  wire multm_reduce_mulsc_mulb_ps97;
  wire multm_reduce_mulsc_mulb_ps98;
  wire multm_reduce_mulsc_mulb_ps99;
  wire multm_reduce_mulsc_mulb_ps100;
  wire multm_reduce_mulsc_mulb_ps101;
  wire multm_reduce_mulsc_mulb_ps102;
  wire multm_reduce_mulsc_mulb_ps103;
  wire multm_reduce_mulsc_mulb_ps104;
  wire multm_reduce_mulsc_mulb_ps105;
  wire multm_reduce_mulsc_mulb_ps106;
  wire multm_reduce_mulsc_mulb_ps107;
  wire multm_reduce_mulsc_mulb_ps108;
  wire multm_reduce_mulsc_mulb_ps109;
  wire multm_reduce_mulsc_mulb_ps110;
  wire multm_reduce_mulsc_mulb_ps111;
  wire multm_reduce_mulsc_mulb_ps112;
  wire multm_reduce_mulsc_mulb_ps113;
  wire multm_reduce_mulsc_mulb_ps114;
  wire multm_reduce_mulsc_mulb_ps115;
  wire multm_reduce_mulsc_mulb_ps116;
  wire multm_reduce_mulsc_mulb_ps117;
  wire multm_reduce_mulsc_mulb_ps118;
  wire multm_reduce_mulsc_mulb_ps119;
  wire multm_reduce_mulsc_mulb_ps120;
  wire multm_reduce_mulsc_mulb_ps121;
  wire multm_reduce_mulsc_mulb_ps122;
  wire multm_reduce_mulsc_mulb_ps123;
  wire multm_reduce_mulsc_mulb_ps124;
  wire multm_reduce_mulsc_mulb_ps125;
  wire multm_reduce_mulsc_mulb_ps126;
  wire multm_reduce_mulsc_mulb_ps127;
  wire multm_reduce_mulsc_mulb_ps128;
  wire multm_reduce_mulsc_mulb_ps129;
  wire multm_reduce_mulsc_mulb_ps130;
  wire multm_reduce_mulsc_mulb_ps131;
  wire multm_reduce_mulsc_mulb_ps132;
  wire multm_reduce_mulsc_mulb_ps133;
  wire multm_reduce_mulsc_mulb_ps134;
  wire multm_reduce_mulsc_mulb_ps135;
  wire multm_reduce_mulsc_mulb_ps136;
  wire multm_reduce_mulsc_mulb_ps137;
  wire multm_reduce_mulsc_mulb_ps138;
  wire multm_reduce_mulsc_mulb_ps139;
  wire multm_reduce_mulsc_mulb_ps140;
  wire multm_reduce_mulsc_mulb_ps141;
  wire multm_reduce_mulsc_mulb_ps142;
  wire multm_reduce_mulsc_mulb_ps143;
  wire multm_reduce_mulsc_mulb_ps144;
  wire multm_reduce_mulsc_mulb_ps145;
  wire multm_reduce_mulsc_mulb_ps146;
  wire multm_reduce_mulsc_mulb_ps147;
  wire multm_reduce_mulsc_mulb_ps148;
  wire multm_reduce_mulsc_mulb_ps149;
  wire multm_reduce_mulsc_mulb_ps150;
  wire multm_reduce_mulsc_mulb_ps151;
  wire multm_reduce_mulsc_mulb_ps152;
  wire multm_reduce_mulsc_mulb_ps153;
  wire multm_reduce_mulsc_mulb_ps154;
  wire multm_reduce_mulsc_mulb_ps155;
  wire multm_reduce_mulsc_mulb_ps156;
  wire multm_reduce_mulsc_mulb_ps157;
  wire multm_reduce_mulsc_mulb_ps158;
  wire multm_reduce_mulsc_mulb_ps159;
  wire multm_reduce_mulsc_mulb_ps160;
  wire multm_reduce_mulsc_mulb_ps161;
  wire multm_reduce_mulsc_mulb_ps162;
  wire multm_reduce_mulsc_mulb_ps163;
  wire multm_reduce_mulsc_mulb_ps164;
  wire multm_reduce_mulsc_mulb_ps165;
  wire multm_reduce_mulsc_mulb_ps166;
  wire multm_reduce_mulsc_mulb_ps167;
  wire multm_reduce_mulsc_mulb_ps168;
  wire multm_reduce_mulsc_mulb_ps169;
  wire multm_reduce_mulsc_mulb_ps170;
  wire multm_reduce_mulsc_mulb_ps171;
  wire multm_reduce_mulsc_mulb_ps172;
  wire multm_reduce_mulsc_mulb_ps173;
  wire multm_reduce_mulsc_mulb_ps174;
  wire multm_reduce_mulsc_mulb_ps175;
  wire multm_reduce_mulsc_mulb_ps176;
  wire multm_reduce_mulsc_mulb_ps177;
  wire multm_reduce_mulsc_mulb_ps178;
  wire multm_reduce_mulsc_mulb_ps179;
  wire multm_reduce_mulsc_mulb_ps180;
  wire multm_reduce_mulsc_mulb_ps181;
  wire multm_reduce_mulsc_mulb_ps182;
  wire multm_reduce_mulsc_mulb_sq0;
  wire multm_reduce_mulsc_mulb_sq1;
  wire multm_reduce_mulsc_mulb_sq2;
  wire multm_reduce_mulsc_mulb_sq3;
  wire multm_reduce_mulsc_mulb_sq4;
  wire multm_reduce_mulsc_mulb_sq5;
  wire multm_reduce_mulsc_mulb_sq6;
  wire multm_reduce_mulsc_mulb_sq7;
  wire multm_reduce_mulsc_mulb_sq8;
  wire multm_reduce_mulsc_mulb_sq9;
  wire multm_reduce_mulsc_mulb_sq10;
  wire multm_reduce_mulsc_mulb_sq11;
  wire multm_reduce_mulsc_mulb_sq12;
  wire multm_reduce_mulsc_mulb_sq13;
  wire multm_reduce_mulsc_mulb_sq14;
  wire multm_reduce_mulsc_mulb_sq15;
  wire multm_reduce_mulsc_mulb_sq16;
  wire multm_reduce_mulsc_mulb_sq17;
  wire multm_reduce_mulsc_mulb_sq18;
  wire multm_reduce_mulsc_mulb_sq19;
  wire multm_reduce_mulsc_mulb_sq20;
  wire multm_reduce_mulsc_mulb_sq21;
  wire multm_reduce_mulsc_mulb_sq22;
  wire multm_reduce_mulsc_mulb_sq23;
  wire multm_reduce_mulsc_mulb_sq24;
  wire multm_reduce_mulsc_mulb_sq25;
  wire multm_reduce_mulsc_mulb_sq26;
  wire multm_reduce_mulsc_mulb_sq27;
  wire multm_reduce_mulsc_mulb_sq28;
  wire multm_reduce_mulsc_mulb_sq29;
  wire multm_reduce_mulsc_mulb_sq30;
  wire multm_reduce_mulsc_mulb_sq31;
  wire multm_reduce_mulsc_mulb_sq32;
  wire multm_reduce_mulsc_mulb_sq33;
  wire multm_reduce_mulsc_mulb_sq34;
  wire multm_reduce_mulsc_mulb_sq35;
  wire multm_reduce_mulsc_mulb_sq36;
  wire multm_reduce_mulsc_mulb_sq37;
  wire multm_reduce_mulsc_mulb_sq38;
  wire multm_reduce_mulsc_mulb_sq39;
  wire multm_reduce_mulsc_mulb_sq40;
  wire multm_reduce_mulsc_mulb_sq41;
  wire multm_reduce_mulsc_mulb_sq42;
  wire multm_reduce_mulsc_mulb_sq43;
  wire multm_reduce_mulsc_mulb_sq44;
  wire multm_reduce_mulsc_mulb_sq45;
  wire multm_reduce_mulsc_mulb_sq46;
  wire multm_reduce_mulsc_mulb_sq47;
  wire multm_reduce_mulsc_mulb_sq48;
  wire multm_reduce_mulsc_mulb_sq49;
  wire multm_reduce_mulsc_mulb_sq50;
  wire multm_reduce_mulsc_mulb_sq51;
  wire multm_reduce_mulsc_mulb_sq52;
  wire multm_reduce_mulsc_mulb_sq53;
  wire multm_reduce_mulsc_mulb_sq54;
  wire multm_reduce_mulsc_mulb_sq55;
  wire multm_reduce_mulsc_mulb_sq56;
  wire multm_reduce_mulsc_mulb_sq57;
  wire multm_reduce_mulsc_mulb_sq58;
  wire multm_reduce_mulsc_mulb_sq59;
  wire multm_reduce_mulsc_mulb_sq60;
  wire multm_reduce_mulsc_mulb_sq61;
  wire multm_reduce_mulsc_mulb_sq62;
  wire multm_reduce_mulsc_mulb_sq63;
  wire multm_reduce_mulsc_mulb_sq64;
  wire multm_reduce_mulsc_mulb_sq65;
  wire multm_reduce_mulsc_mulb_sq66;
  wire multm_reduce_mulsc_mulb_sq67;
  wire multm_reduce_mulsc_mulb_sq68;
  wire multm_reduce_mulsc_mulb_sq69;
  wire multm_reduce_mulsc_mulb_sq70;
  wire multm_reduce_mulsc_mulb_sq71;
  wire multm_reduce_mulsc_mulb_sq72;
  wire multm_reduce_mulsc_mulb_sq73;
  wire multm_reduce_mulsc_mulb_sq74;
  wire multm_reduce_mulsc_mulb_sq75;
  wire multm_reduce_mulsc_mulb_sq76;
  wire multm_reduce_mulsc_mulb_sq77;
  wire multm_reduce_mulsc_mulb_sq78;
  wire multm_reduce_mulsc_mulb_sq79;
  wire multm_reduce_mulsc_mulb_sq80;
  wire multm_reduce_mulsc_mulb_sq81;
  wire multm_reduce_mulsc_mulb_sq82;
  wire multm_reduce_mulsc_mulb_sq83;
  wire multm_reduce_mulsc_mulb_sq84;
  wire multm_reduce_mulsc_mulb_sq85;
  wire multm_reduce_mulsc_mulb_sq86;
  wire multm_reduce_mulsc_mulb_sq87;
  wire multm_reduce_mulsc_mulb_sq88;
  wire multm_reduce_mulsc_mulb_sq89;
  wire multm_reduce_mulsc_mulb_sq90;
  wire multm_reduce_mulsc_mulb_sq91;
  wire multm_reduce_mulsc_mulb_sq92;
  wire multm_reduce_mulsc_mulb_sq93;
  wire multm_reduce_mulsc_mulb_sq94;
  wire multm_reduce_mulsc_mulb_sq95;
  wire multm_reduce_mulsc_mulb_sq96;
  wire multm_reduce_mulsc_mulb_sq97;
  wire multm_reduce_mulsc_mulb_sq98;
  wire multm_reduce_mulsc_mulb_sq99;
  wire multm_reduce_mulsc_mulb_sq100;
  wire multm_reduce_mulsc_mulb_sq101;
  wire multm_reduce_mulsc_mulb_sq102;
  wire multm_reduce_mulsc_mulb_sq103;
  wire multm_reduce_mulsc_mulb_sq104;
  wire multm_reduce_mulsc_mulb_sq105;
  wire multm_reduce_mulsc_mulb_sq106;
  wire multm_reduce_mulsc_mulb_sq107;
  wire multm_reduce_mulsc_mulb_sq108;
  wire multm_reduce_mulsc_mulb_sq109;
  wire multm_reduce_mulsc_mulb_sq110;
  wire multm_reduce_mulsc_mulb_sq111;
  wire multm_reduce_mulsc_mulb_sq112;
  wire multm_reduce_mulsc_mulb_sq113;
  wire multm_reduce_mulsc_mulb_sq114;
  wire multm_reduce_mulsc_mulb_sq115;
  wire multm_reduce_mulsc_mulb_sq116;
  wire multm_reduce_mulsc_mulb_sq117;
  wire multm_reduce_mulsc_mulb_sq118;
  wire multm_reduce_mulsc_mulb_sq119;
  wire multm_reduce_mulsc_mulb_sq120;
  wire multm_reduce_mulsc_mulb_sq121;
  wire multm_reduce_mulsc_mulb_sq122;
  wire multm_reduce_mulsc_mulb_sq123;
  wire multm_reduce_mulsc_mulb_sq124;
  wire multm_reduce_mulsc_mulb_sq125;
  wire multm_reduce_mulsc_mulb_sq126;
  wire multm_reduce_mulsc_mulb_sq127;
  wire multm_reduce_mulsc_mulb_sq128;
  wire multm_reduce_mulsc_mulb_sq129;
  wire multm_reduce_mulsc_mulb_sq130;
  wire multm_reduce_mulsc_mulb_sq131;
  wire multm_reduce_mulsc_mulb_sq132;
  wire multm_reduce_mulsc_mulb_sq133;
  wire multm_reduce_mulsc_mulb_sq134;
  wire multm_reduce_mulsc_mulb_sq135;
  wire multm_reduce_mulsc_mulb_sq136;
  wire multm_reduce_mulsc_mulb_sq137;
  wire multm_reduce_mulsc_mulb_sq138;
  wire multm_reduce_mulsc_mulb_sq139;
  wire multm_reduce_mulsc_mulb_sq140;
  wire multm_reduce_mulsc_mulb_sq141;
  wire multm_reduce_mulsc_mulb_sq142;
  wire multm_reduce_mulsc_mulb_sq143;
  wire multm_reduce_mulsc_mulb_sq144;
  wire multm_reduce_mulsc_mulb_sq145;
  wire multm_reduce_mulsc_mulb_sq146;
  wire multm_reduce_mulsc_mulb_sq147;
  wire multm_reduce_mulsc_mulb_sq148;
  wire multm_reduce_mulsc_mulb_sq149;
  wire multm_reduce_mulsc_mulb_sq150;
  wire multm_reduce_mulsc_mulb_sq151;
  wire multm_reduce_mulsc_mulb_sq152;
  wire multm_reduce_mulsc_mulb_sq153;
  wire multm_reduce_mulsc_mulb_sq154;
  wire multm_reduce_mulsc_mulb_sq155;
  wire multm_reduce_mulsc_mulb_sq156;
  wire multm_reduce_mulsc_mulb_sq157;
  wire multm_reduce_mulsc_mulb_sq158;
  wire multm_reduce_mulsc_mulb_sq159;
  wire multm_reduce_mulsc_mulb_sq160;
  wire multm_reduce_mulsc_mulb_sq161;
  wire multm_reduce_mulsc_mulb_sq162;
  wire multm_reduce_mulsc_mulb_sq163;
  wire multm_reduce_mulsc_mulb_sq164;
  wire multm_reduce_mulsc_mulb_sq165;
  wire multm_reduce_mulsc_mulb_sq166;
  wire multm_reduce_mulsc_mulb_sq167;
  wire multm_reduce_mulsc_mulb_sq168;
  wire multm_reduce_mulsc_mulb_sq169;
  wire multm_reduce_mulsc_mulb_sq170;
  wire multm_reduce_mulsc_mulb_sq171;
  wire multm_reduce_mulsc_mulb_sq172;
  wire multm_reduce_mulsc_mulb_sq173;
  wire multm_reduce_mulsc_mulb_sq174;
  wire multm_reduce_mulsc_mulb_sq175;
  wire multm_reduce_mulsc_mulb_sq176;
  wire multm_reduce_mulsc_mulb_sq177;
  wire multm_reduce_mulsc_mulb_sq178;
  wire multm_reduce_mulsc_mulb_sq179;
  wire multm_reduce_mulsc_mulb_sq180;
  wire multm_reduce_mulsc_mulb_sq181;
  wire multm_reduce_mulsc_mulb_sq182;
  wire multm_reduce_mulsc_mulb_sq183;
  wire multm_reduce_mulsc_mulb_yoc0;
  wire multm_reduce_mulsc_mulb_yoc1;
  wire multm_reduce_mulsc_mulb_yoc2;
  wire multm_reduce_mulsc_mulb_yoc3;
  wire multm_reduce_mulsc_mulb_yoc4;
  wire multm_reduce_mulsc_mulb_yoc5;
  wire multm_reduce_mulsc_mulb_yoc6;
  wire multm_reduce_mulsc_mulb_yoc7;
  wire multm_reduce_mulsc_mulb_yoc8;
  wire multm_reduce_mulsc_mulb_yoc9;
  wire multm_reduce_mulsc_mulb_yoc10;
  wire multm_reduce_mulsc_mulb_yoc11;
  wire multm_reduce_mulsc_mulb_yoc12;
  wire multm_reduce_mulsc_mulb_yoc13;
  wire multm_reduce_mulsc_mulb_yoc14;
  wire multm_reduce_mulsc_mulb_yoc15;
  wire multm_reduce_mulsc_mulb_yoc16;
  wire multm_reduce_mulsc_mulb_yoc17;
  wire multm_reduce_mulsc_mulb_yoc18;
  wire multm_reduce_mulsc_mulb_yoc19;
  wire multm_reduce_mulsc_mulb_yoc20;
  wire multm_reduce_mulsc_mulb_yoc21;
  wire multm_reduce_mulsc_mulb_yoc22;
  wire multm_reduce_mulsc_mulb_yoc23;
  wire multm_reduce_mulsc_mulb_yoc24;
  wire multm_reduce_mulsc_mulb_yoc25;
  wire multm_reduce_mulsc_mulb_yoc26;
  wire multm_reduce_mulsc_mulb_yoc27;
  wire multm_reduce_mulsc_mulb_yoc28;
  wire multm_reduce_mulsc_mulb_yoc29;
  wire multm_reduce_mulsc_mulb_yoc30;
  wire multm_reduce_mulsc_mulb_yoc31;
  wire multm_reduce_mulsc_mulb_yoc32;
  wire multm_reduce_mulsc_mulb_yoc33;
  wire multm_reduce_mulsc_mulb_yoc34;
  wire multm_reduce_mulsc_mulb_yoc35;
  wire multm_reduce_mulsc_mulb_yoc36;
  wire multm_reduce_mulsc_mulb_yoc37;
  wire multm_reduce_mulsc_mulb_yoc38;
  wire multm_reduce_mulsc_mulb_yoc39;
  wire multm_reduce_mulsc_mulb_yoc40;
  wire multm_reduce_mulsc_mulb_yoc41;
  wire multm_reduce_mulsc_mulb_yoc42;
  wire multm_reduce_mulsc_mulb_yoc43;
  wire multm_reduce_mulsc_mulb_yoc44;
  wire multm_reduce_mulsc_mulb_yoc45;
  wire multm_reduce_mulsc_mulb_yoc46;
  wire multm_reduce_mulsc_mulb_yoc47;
  wire multm_reduce_mulsc_mulb_yoc48;
  wire multm_reduce_mulsc_mulb_yoc49;
  wire multm_reduce_mulsc_mulb_yoc50;
  wire multm_reduce_mulsc_mulb_yoc51;
  wire multm_reduce_mulsc_mulb_yoc52;
  wire multm_reduce_mulsc_mulb_yoc53;
  wire multm_reduce_mulsc_mulb_yoc54;
  wire multm_reduce_mulsc_mulb_yoc55;
  wire multm_reduce_mulsc_mulb_yoc56;
  wire multm_reduce_mulsc_mulb_yoc57;
  wire multm_reduce_mulsc_mulb_yoc58;
  wire multm_reduce_mulsc_mulb_yoc59;
  wire multm_reduce_mulsc_mulb_yoc60;
  wire multm_reduce_mulsc_mulb_yoc61;
  wire multm_reduce_mulsc_mulb_yoc62;
  wire multm_reduce_mulsc_mulb_yoc63;
  wire multm_reduce_mulsc_mulb_yoc64;
  wire multm_reduce_mulsc_mulb_yoc65;
  wire multm_reduce_mulsc_mulb_yoc66;
  wire multm_reduce_mulsc_mulb_yoc67;
  wire multm_reduce_mulsc_mulb_yoc68;
  wire multm_reduce_mulsc_mulb_yoc69;
  wire multm_reduce_mulsc_mulb_yoc70;
  wire multm_reduce_mulsc_mulb_yoc71;
  wire multm_reduce_mulsc_mulb_yoc72;
  wire multm_reduce_mulsc_mulb_yoc73;
  wire multm_reduce_mulsc_mulb_yoc74;
  wire multm_reduce_mulsc_mulb_yoc75;
  wire multm_reduce_mulsc_mulb_yoc76;
  wire multm_reduce_mulsc_mulb_yoc77;
  wire multm_reduce_mulsc_mulb_yoc78;
  wire multm_reduce_mulsc_mulb_yoc79;
  wire multm_reduce_mulsc_mulb_yoc80;
  wire multm_reduce_mulsc_mulb_yoc81;
  wire multm_reduce_mulsc_mulb_yoc82;
  wire multm_reduce_mulsc_mulb_yoc83;
  wire multm_reduce_mulsc_mulb_yoc84;
  wire multm_reduce_mulsc_mulb_yoc85;
  wire multm_reduce_mulsc_mulb_yoc86;
  wire multm_reduce_mulsc_mulb_yoc87;
  wire multm_reduce_mulsc_mulb_yoc88;
  wire multm_reduce_mulsc_mulb_yoc89;
  wire multm_reduce_mulsc_mulb_yoc90;
  wire multm_reduce_mulsc_mulb_yoc91;
  wire multm_reduce_mulsc_mulb_yoc92;
  wire multm_reduce_mulsc_mulb_yoc93;
  wire multm_reduce_mulsc_mulb_yoc94;
  wire multm_reduce_mulsc_mulb_yoc95;
  wire multm_reduce_mulsc_mulb_yoc96;
  wire multm_reduce_mulsc_mulb_yoc97;
  wire multm_reduce_mulsc_mulb_yoc98;
  wire multm_reduce_mulsc_mulb_yoc99;
  wire multm_reduce_mulsc_mulb_yoc100;
  wire multm_reduce_mulsc_mulb_yoc101;
  wire multm_reduce_mulsc_mulb_yoc102;
  wire multm_reduce_mulsc_mulb_yoc103;
  wire multm_reduce_mulsc_mulb_yoc104;
  wire multm_reduce_mulsc_mulb_yoc105;
  wire multm_reduce_mulsc_mulb_yoc106;
  wire multm_reduce_mulsc_mulb_yoc107;
  wire multm_reduce_mulsc_mulb_yoc108;
  wire multm_reduce_mulsc_mulb_yoc109;
  wire multm_reduce_mulsc_mulb_yoc110;
  wire multm_reduce_mulsc_mulb_yoc111;
  wire multm_reduce_mulsc_mulb_yoc112;
  wire multm_reduce_mulsc_mulb_yoc113;
  wire multm_reduce_mulsc_mulb_yoc114;
  wire multm_reduce_mulsc_mulb_yoc115;
  wire multm_reduce_mulsc_mulb_yoc116;
  wire multm_reduce_mulsc_mulb_yoc117;
  wire multm_reduce_mulsc_mulb_yoc118;
  wire multm_reduce_mulsc_mulb_yoc119;
  wire multm_reduce_mulsc_mulb_yoc120;
  wire multm_reduce_mulsc_mulb_yoc121;
  wire multm_reduce_mulsc_mulb_yoc122;
  wire multm_reduce_mulsc_mulb_yoc123;
  wire multm_reduce_mulsc_mulb_yoc124;
  wire multm_reduce_mulsc_mulb_yoc125;
  wire multm_reduce_mulsc_mulb_yoc126;
  wire multm_reduce_mulsc_mulb_yoc127;
  wire multm_reduce_mulsc_mulb_yoc128;
  wire multm_reduce_mulsc_mulb_yoc129;
  wire multm_reduce_mulsc_mulb_yoc130;
  wire multm_reduce_mulsc_mulb_yoc131;
  wire multm_reduce_mulsc_mulb_yoc132;
  wire multm_reduce_mulsc_mulb_yoc133;
  wire multm_reduce_mulsc_mulb_yoc134;
  wire multm_reduce_mulsc_mulb_yoc135;
  wire multm_reduce_mulsc_mulb_yoc136;
  wire multm_reduce_mulsc_mulb_yoc137;
  wire multm_reduce_mulsc_mulb_yoc138;
  wire multm_reduce_mulsc_mulb_yoc139;
  wire multm_reduce_mulsc_mulb_yoc140;
  wire multm_reduce_mulsc_mulb_yoc141;
  wire multm_reduce_mulsc_mulb_yoc142;
  wire multm_reduce_mulsc_mulb_yoc143;
  wire multm_reduce_mulsc_mulb_yoc144;
  wire multm_reduce_mulsc_mulb_yoc145;
  wire multm_reduce_mulsc_mulb_yoc146;
  wire multm_reduce_mulsc_mulb_yoc147;
  wire multm_reduce_mulsc_mulb_yoc148;
  wire multm_reduce_mulsc_mulb_yoc149;
  wire multm_reduce_mulsc_mulb_yoc150;
  wire multm_reduce_mulsc_mulb_yoc151;
  wire multm_reduce_mulsc_mulb_yoc152;
  wire multm_reduce_mulsc_mulb_yoc153;
  wire multm_reduce_mulsc_mulb_yoc154;
  wire multm_reduce_mulsc_mulb_yoc155;
  wire multm_reduce_mulsc_mulb_yoc156;
  wire multm_reduce_mulsc_mulb_yoc157;
  wire multm_reduce_mulsc_mulb_yoc158;
  wire multm_reduce_mulsc_mulb_yoc159;
  wire multm_reduce_mulsc_mulb_yoc160;
  wire multm_reduce_mulsc_mulb_yoc161;
  wire multm_reduce_mulsc_mulb_yoc162;
  wire multm_reduce_mulsc_mulb_yoc163;
  wire multm_reduce_mulsc_mulb_yoc164;
  wire multm_reduce_mulsc_mulb_yoc165;
  wire multm_reduce_mulsc_mulb_yoc166;
  wire multm_reduce_mulsc_mulb_yoc167;
  wire multm_reduce_mulsc_mulb_yoc168;
  wire multm_reduce_mulsc_mulb_yoc169;
  wire multm_reduce_mulsc_mulb_yoc170;
  wire multm_reduce_mulsc_mulb_yoc171;
  wire multm_reduce_mulsc_mulb_yoc172;
  wire multm_reduce_mulsc_mulb_yoc173;
  wire multm_reduce_mulsc_mulb_yoc174;
  wire multm_reduce_mulsc_mulb_yoc175;
  wire multm_reduce_mulsc_mulb_yoc176;
  wire multm_reduce_mulsc_mulb_yoc177;
  wire multm_reduce_mulsc_mulb_yoc178;
  wire multm_reduce_mulsc_mulb_yoc179;
  wire multm_reduce_mulsc_mulb_yoc180;
  wire multm_reduce_mulsc_mulb_yoc181;
  wire multm_reduce_mulsc_mulb_yoc182;
  wire multm_reduce_mulsc_mulb_yoc183;
  wire multm_reduce_mulsc_mulb_yos0;
  wire multm_reduce_mulsc_mulb_yos1;
  wire multm_reduce_mulsc_mulb_yos2;
  wire multm_reduce_mulsc_mulb_yos3;
  wire multm_reduce_mulsc_mulb_yos4;
  wire multm_reduce_mulsc_mulb_yos5;
  wire multm_reduce_mulsc_mulb_yos6;
  wire multm_reduce_mulsc_mulb_yos7;
  wire multm_reduce_mulsc_mulb_yos8;
  wire multm_reduce_mulsc_mulb_yos9;
  wire multm_reduce_mulsc_mulb_yos10;
  wire multm_reduce_mulsc_mulb_yos11;
  wire multm_reduce_mulsc_mulb_yos12;
  wire multm_reduce_mulsc_mulb_yos13;
  wire multm_reduce_mulsc_mulb_yos14;
  wire multm_reduce_mulsc_mulb_yos15;
  wire multm_reduce_mulsc_mulb_yos16;
  wire multm_reduce_mulsc_mulb_yos17;
  wire multm_reduce_mulsc_mulb_yos18;
  wire multm_reduce_mulsc_mulb_yos19;
  wire multm_reduce_mulsc_mulb_yos20;
  wire multm_reduce_mulsc_mulb_yos21;
  wire multm_reduce_mulsc_mulb_yos22;
  wire multm_reduce_mulsc_mulb_yos23;
  wire multm_reduce_mulsc_mulb_yos24;
  wire multm_reduce_mulsc_mulb_yos25;
  wire multm_reduce_mulsc_mulb_yos26;
  wire multm_reduce_mulsc_mulb_yos27;
  wire multm_reduce_mulsc_mulb_yos28;
  wire multm_reduce_mulsc_mulb_yos29;
  wire multm_reduce_mulsc_mulb_yos30;
  wire multm_reduce_mulsc_mulb_yos31;
  wire multm_reduce_mulsc_mulb_yos32;
  wire multm_reduce_mulsc_mulb_yos33;
  wire multm_reduce_mulsc_mulb_yos34;
  wire multm_reduce_mulsc_mulb_yos35;
  wire multm_reduce_mulsc_mulb_yos36;
  wire multm_reduce_mulsc_mulb_yos37;
  wire multm_reduce_mulsc_mulb_yos38;
  wire multm_reduce_mulsc_mulb_yos39;
  wire multm_reduce_mulsc_mulb_yos40;
  wire multm_reduce_mulsc_mulb_yos41;
  wire multm_reduce_mulsc_mulb_yos42;
  wire multm_reduce_mulsc_mulb_yos43;
  wire multm_reduce_mulsc_mulb_yos44;
  wire multm_reduce_mulsc_mulb_yos45;
  wire multm_reduce_mulsc_mulb_yos46;
  wire multm_reduce_mulsc_mulb_yos47;
  wire multm_reduce_mulsc_mulb_yos48;
  wire multm_reduce_mulsc_mulb_yos49;
  wire multm_reduce_mulsc_mulb_yos50;
  wire multm_reduce_mulsc_mulb_yos51;
  wire multm_reduce_mulsc_mulb_yos52;
  wire multm_reduce_mulsc_mulb_yos53;
  wire multm_reduce_mulsc_mulb_yos54;
  wire multm_reduce_mulsc_mulb_yos55;
  wire multm_reduce_mulsc_mulb_yos56;
  wire multm_reduce_mulsc_mulb_yos57;
  wire multm_reduce_mulsc_mulb_yos58;
  wire multm_reduce_mulsc_mulb_yos59;
  wire multm_reduce_mulsc_mulb_yos60;
  wire multm_reduce_mulsc_mulb_yos61;
  wire multm_reduce_mulsc_mulb_yos62;
  wire multm_reduce_mulsc_mulb_yos63;
  wire multm_reduce_mulsc_mulb_yos64;
  wire multm_reduce_mulsc_mulb_yos65;
  wire multm_reduce_mulsc_mulb_yos66;
  wire multm_reduce_mulsc_mulb_yos67;
  wire multm_reduce_mulsc_mulb_yos68;
  wire multm_reduce_mulsc_mulb_yos69;
  wire multm_reduce_mulsc_mulb_yos70;
  wire multm_reduce_mulsc_mulb_yos71;
  wire multm_reduce_mulsc_mulb_yos72;
  wire multm_reduce_mulsc_mulb_yos73;
  wire multm_reduce_mulsc_mulb_yos74;
  wire multm_reduce_mulsc_mulb_yos75;
  wire multm_reduce_mulsc_mulb_yos76;
  wire multm_reduce_mulsc_mulb_yos77;
  wire multm_reduce_mulsc_mulb_yos78;
  wire multm_reduce_mulsc_mulb_yos79;
  wire multm_reduce_mulsc_mulb_yos80;
  wire multm_reduce_mulsc_mulb_yos81;
  wire multm_reduce_mulsc_mulb_yos82;
  wire multm_reduce_mulsc_mulb_yos83;
  wire multm_reduce_mulsc_mulb_yos84;
  wire multm_reduce_mulsc_mulb_yos85;
  wire multm_reduce_mulsc_mulb_yos86;
  wire multm_reduce_mulsc_mulb_yos87;
  wire multm_reduce_mulsc_mulb_yos88;
  wire multm_reduce_mulsc_mulb_yos89;
  wire multm_reduce_mulsc_mulb_yos90;
  wire multm_reduce_mulsc_mulb_yos91;
  wire multm_reduce_mulsc_mulb_yos92;
  wire multm_reduce_mulsc_mulb_yos93;
  wire multm_reduce_mulsc_mulb_yos94;
  wire multm_reduce_mulsc_mulb_yos95;
  wire multm_reduce_mulsc_mulb_yos96;
  wire multm_reduce_mulsc_mulb_yos97;
  wire multm_reduce_mulsc_mulb_yos98;
  wire multm_reduce_mulsc_mulb_yos99;
  wire multm_reduce_mulsc_mulb_yos100;
  wire multm_reduce_mulsc_mulb_yos101;
  wire multm_reduce_mulsc_mulb_yos102;
  wire multm_reduce_mulsc_mulb_yos103;
  wire multm_reduce_mulsc_mulb_yos104;
  wire multm_reduce_mulsc_mulb_yos105;
  wire multm_reduce_mulsc_mulb_yos106;
  wire multm_reduce_mulsc_mulb_yos107;
  wire multm_reduce_mulsc_mulb_yos108;
  wire multm_reduce_mulsc_mulb_yos109;
  wire multm_reduce_mulsc_mulb_yos110;
  wire multm_reduce_mulsc_mulb_yos111;
  wire multm_reduce_mulsc_mulb_yos112;
  wire multm_reduce_mulsc_mulb_yos113;
  wire multm_reduce_mulsc_mulb_yos114;
  wire multm_reduce_mulsc_mulb_yos115;
  wire multm_reduce_mulsc_mulb_yos116;
  wire multm_reduce_mulsc_mulb_yos117;
  wire multm_reduce_mulsc_mulb_yos118;
  wire multm_reduce_mulsc_mulb_yos119;
  wire multm_reduce_mulsc_mulb_yos120;
  wire multm_reduce_mulsc_mulb_yos121;
  wire multm_reduce_mulsc_mulb_yos122;
  wire multm_reduce_mulsc_mulb_yos123;
  wire multm_reduce_mulsc_mulb_yos124;
  wire multm_reduce_mulsc_mulb_yos125;
  wire multm_reduce_mulsc_mulb_yos126;
  wire multm_reduce_mulsc_mulb_yos127;
  wire multm_reduce_mulsc_mulb_yos128;
  wire multm_reduce_mulsc_mulb_yos129;
  wire multm_reduce_mulsc_mulb_yos130;
  wire multm_reduce_mulsc_mulb_yos131;
  wire multm_reduce_mulsc_mulb_yos132;
  wire multm_reduce_mulsc_mulb_yos133;
  wire multm_reduce_mulsc_mulb_yos134;
  wire multm_reduce_mulsc_mulb_yos135;
  wire multm_reduce_mulsc_mulb_yos136;
  wire multm_reduce_mulsc_mulb_yos137;
  wire multm_reduce_mulsc_mulb_yos138;
  wire multm_reduce_mulsc_mulb_yos139;
  wire multm_reduce_mulsc_mulb_yos140;
  wire multm_reduce_mulsc_mulb_yos141;
  wire multm_reduce_mulsc_mulb_yos142;
  wire multm_reduce_mulsc_mulb_yos143;
  wire multm_reduce_mulsc_mulb_yos144;
  wire multm_reduce_mulsc_mulb_yos145;
  wire multm_reduce_mulsc_mulb_yos146;
  wire multm_reduce_mulsc_mulb_yos147;
  wire multm_reduce_mulsc_mulb_yos148;
  wire multm_reduce_mulsc_mulb_yos149;
  wire multm_reduce_mulsc_mulb_yos150;
  wire multm_reduce_mulsc_mulb_yos151;
  wire multm_reduce_mulsc_mulb_yos152;
  wire multm_reduce_mulsc_mulb_yos153;
  wire multm_reduce_mulsc_mulb_yos154;
  wire multm_reduce_mulsc_mulb_yos155;
  wire multm_reduce_mulsc_mulb_yos156;
  wire multm_reduce_mulsc_mulb_yos157;
  wire multm_reduce_mulsc_mulb_yos158;
  wire multm_reduce_mulsc_mulb_yos159;
  wire multm_reduce_mulsc_mulb_yos160;
  wire multm_reduce_mulsc_mulb_yos161;
  wire multm_reduce_mulsc_mulb_yos162;
  wire multm_reduce_mulsc_mulb_yos163;
  wire multm_reduce_mulsc_mulb_yos164;
  wire multm_reduce_mulsc_mulb_yos165;
  wire multm_reduce_mulsc_mulb_yos166;
  wire multm_reduce_mulsc_mulb_yos167;
  wire multm_reduce_mulsc_mulb_yos168;
  wire multm_reduce_mulsc_mulb_yos169;
  wire multm_reduce_mulsc_mulb_yos170;
  wire multm_reduce_mulsc_mulb_yos171;
  wire multm_reduce_mulsc_mulb_yos172;
  wire multm_reduce_mulsc_mulb_yos173;
  wire multm_reduce_mulsc_mulb_yos174;
  wire multm_reduce_mulsc_mulb_yos175;
  wire multm_reduce_mulsc_mulb_yos176;
  wire multm_reduce_mulsc_mulb_yos177;
  wire multm_reduce_mulsc_mulb_yos178;
  wire multm_reduce_mulsc_mulb_yos179;
  wire multm_reduce_mulsc_mulb_yos180;
  wire multm_reduce_mulsc_mulb_yos181;
  wire multm_reduce_mulsc_mulb_yos182;
  wire multm_reduce_mulsc_mulb_yos183;
  wire multm_reduce_mulsc_shrsc_cq0;
  wire multm_reduce_mulsc_shrsc_cq1;
  wire multm_reduce_mulsc_shrsc_cq2;
  wire multm_reduce_mulsc_shrsc_cq3;
  wire multm_reduce_mulsc_shrsc_cq4;
  wire multm_reduce_mulsc_shrsc_cq5;
  wire multm_reduce_mulsc_shrsc_cq6;
  wire multm_reduce_mulsc_shrsc_cq7;
  wire multm_reduce_mulsc_shrsc_cq8;
  wire multm_reduce_mulsc_shrsc_cq9;
  wire multm_reduce_mulsc_shrsc_cq10;
  wire multm_reduce_mulsc_shrsc_cq11;
  wire multm_reduce_mulsc_shrsc_cq12;
  wire multm_reduce_mulsc_shrsc_cq13;
  wire multm_reduce_mulsc_shrsc_cq14;
  wire multm_reduce_mulsc_shrsc_cq15;
  wire multm_reduce_mulsc_shrsc_cq16;
  wire multm_reduce_mulsc_shrsc_cq17;
  wire multm_reduce_mulsc_shrsc_cq18;
  wire multm_reduce_mulsc_shrsc_cq19;
  wire multm_reduce_mulsc_shrsc_cq20;
  wire multm_reduce_mulsc_shrsc_cq21;
  wire multm_reduce_mulsc_shrsc_cq22;
  wire multm_reduce_mulsc_shrsc_cq23;
  wire multm_reduce_mulsc_shrsc_cq24;
  wire multm_reduce_mulsc_shrsc_cq25;
  wire multm_reduce_mulsc_shrsc_cq26;
  wire multm_reduce_mulsc_shrsc_cq27;
  wire multm_reduce_mulsc_shrsc_cq28;
  wire multm_reduce_mulsc_shrsc_cq29;
  wire multm_reduce_mulsc_shrsc_cq30;
  wire multm_reduce_mulsc_shrsc_cq31;
  wire multm_reduce_mulsc_shrsc_cq32;
  wire multm_reduce_mulsc_shrsc_cq33;
  wire multm_reduce_mulsc_shrsc_cq34;
  wire multm_reduce_mulsc_shrsc_cq35;
  wire multm_reduce_mulsc_shrsc_cq36;
  wire multm_reduce_mulsc_shrsc_cq37;
  wire multm_reduce_mulsc_shrsc_cq38;
  wire multm_reduce_mulsc_shrsc_cq39;
  wire multm_reduce_mulsc_shrsc_cq40;
  wire multm_reduce_mulsc_shrsc_cq41;
  wire multm_reduce_mulsc_shrsc_cq42;
  wire multm_reduce_mulsc_shrsc_cq43;
  wire multm_reduce_mulsc_shrsc_cq44;
  wire multm_reduce_mulsc_shrsc_cq45;
  wire multm_reduce_mulsc_shrsc_cq46;
  wire multm_reduce_mulsc_shrsc_cq47;
  wire multm_reduce_mulsc_shrsc_cq48;
  wire multm_reduce_mulsc_shrsc_cq49;
  wire multm_reduce_mulsc_shrsc_cq50;
  wire multm_reduce_mulsc_shrsc_cq51;
  wire multm_reduce_mulsc_shrsc_cq52;
  wire multm_reduce_mulsc_shrsc_cq53;
  wire multm_reduce_mulsc_shrsc_cq54;
  wire multm_reduce_mulsc_shrsc_cq55;
  wire multm_reduce_mulsc_shrsc_cq56;
  wire multm_reduce_mulsc_shrsc_cq57;
  wire multm_reduce_mulsc_shrsc_cq58;
  wire multm_reduce_mulsc_shrsc_cq59;
  wire multm_reduce_mulsc_shrsc_cq60;
  wire multm_reduce_mulsc_shrsc_cq61;
  wire multm_reduce_mulsc_shrsc_cq62;
  wire multm_reduce_mulsc_shrsc_cq63;
  wire multm_reduce_mulsc_shrsc_cq64;
  wire multm_reduce_mulsc_shrsc_cq65;
  wire multm_reduce_mulsc_shrsc_cq66;
  wire multm_reduce_mulsc_shrsc_cq67;
  wire multm_reduce_mulsc_shrsc_cq68;
  wire multm_reduce_mulsc_shrsc_cq69;
  wire multm_reduce_mulsc_shrsc_cq70;
  wire multm_reduce_mulsc_shrsc_cq71;
  wire multm_reduce_mulsc_shrsc_cq72;
  wire multm_reduce_mulsc_shrsc_cq73;
  wire multm_reduce_mulsc_shrsc_cq74;
  wire multm_reduce_mulsc_shrsc_cq75;
  wire multm_reduce_mulsc_shrsc_cq76;
  wire multm_reduce_mulsc_shrsc_cq77;
  wire multm_reduce_mulsc_shrsc_cq78;
  wire multm_reduce_mulsc_shrsc_cq79;
  wire multm_reduce_mulsc_shrsc_cq80;
  wire multm_reduce_mulsc_shrsc_cq81;
  wire multm_reduce_mulsc_shrsc_cq82;
  wire multm_reduce_mulsc_shrsc_cq83;
  wire multm_reduce_mulsc_shrsc_cq84;
  wire multm_reduce_mulsc_shrsc_cq85;
  wire multm_reduce_mulsc_shrsc_cq86;
  wire multm_reduce_mulsc_shrsc_cq87;
  wire multm_reduce_mulsc_shrsc_cq88;
  wire multm_reduce_mulsc_shrsc_cq89;
  wire multm_reduce_mulsc_shrsc_cq90;
  wire multm_reduce_mulsc_shrsc_cq91;
  wire multm_reduce_mulsc_shrsc_cq92;
  wire multm_reduce_mulsc_shrsc_cq93;
  wire multm_reduce_mulsc_shrsc_cq94;
  wire multm_reduce_mulsc_shrsc_cq95;
  wire multm_reduce_mulsc_shrsc_cq96;
  wire multm_reduce_mulsc_shrsc_cq97;
  wire multm_reduce_mulsc_shrsc_cq98;
  wire multm_reduce_mulsc_shrsc_cq99;
  wire multm_reduce_mulsc_shrsc_cq100;
  wire multm_reduce_mulsc_shrsc_cq101;
  wire multm_reduce_mulsc_shrsc_cq102;
  wire multm_reduce_mulsc_shrsc_cq103;
  wire multm_reduce_mulsc_shrsc_cq104;
  wire multm_reduce_mulsc_shrsc_cq105;
  wire multm_reduce_mulsc_shrsc_cq106;
  wire multm_reduce_mulsc_shrsc_cq107;
  wire multm_reduce_mulsc_shrsc_cq108;
  wire multm_reduce_mulsc_shrsc_cq109;
  wire multm_reduce_mulsc_shrsc_cq110;
  wire multm_reduce_mulsc_shrsc_cq111;
  wire multm_reduce_mulsc_shrsc_cq112;
  wire multm_reduce_mulsc_shrsc_cq113;
  wire multm_reduce_mulsc_shrsc_cq114;
  wire multm_reduce_mulsc_shrsc_cq115;
  wire multm_reduce_mulsc_shrsc_cq116;
  wire multm_reduce_mulsc_shrsc_cq117;
  wire multm_reduce_mulsc_shrsc_cq118;
  wire multm_reduce_mulsc_shrsc_cq119;
  wire multm_reduce_mulsc_shrsc_cq120;
  wire multm_reduce_mulsc_shrsc_cq121;
  wire multm_reduce_mulsc_shrsc_cq122;
  wire multm_reduce_mulsc_shrsc_cq123;
  wire multm_reduce_mulsc_shrsc_cq124;
  wire multm_reduce_mulsc_shrsc_cq125;
  wire multm_reduce_mulsc_shrsc_cq126;
  wire multm_reduce_mulsc_shrsc_cq127;
  wire multm_reduce_mulsc_shrsc_cq128;
  wire multm_reduce_mulsc_shrsc_cq129;
  wire multm_reduce_mulsc_shrsc_cq130;
  wire multm_reduce_mulsc_shrsc_cq131;
  wire multm_reduce_mulsc_shrsc_cq132;
  wire multm_reduce_mulsc_shrsc_cq133;
  wire multm_reduce_mulsc_shrsc_cq134;
  wire multm_reduce_mulsc_shrsc_cq135;
  wire multm_reduce_mulsc_shrsc_cq136;
  wire multm_reduce_mulsc_shrsc_cq137;
  wire multm_reduce_mulsc_shrsc_cq138;
  wire multm_reduce_mulsc_shrsc_cq139;
  wire multm_reduce_mulsc_shrsc_cq140;
  wire multm_reduce_mulsc_shrsc_cq141;
  wire multm_reduce_mulsc_shrsc_cq142;
  wire multm_reduce_mulsc_shrsc_cq143;
  wire multm_reduce_mulsc_shrsc_cq144;
  wire multm_reduce_mulsc_shrsc_cq145;
  wire multm_reduce_mulsc_shrsc_cq146;
  wire multm_reduce_mulsc_shrsc_cq147;
  wire multm_reduce_mulsc_shrsc_cq148;
  wire multm_reduce_mulsc_shrsc_cq149;
  wire multm_reduce_mulsc_shrsc_cq150;
  wire multm_reduce_mulsc_shrsc_cq151;
  wire multm_reduce_mulsc_shrsc_cq152;
  wire multm_reduce_mulsc_shrsc_cq153;
  wire multm_reduce_mulsc_shrsc_cq154;
  wire multm_reduce_mulsc_shrsc_cq155;
  wire multm_reduce_mulsc_shrsc_cq156;
  wire multm_reduce_mulsc_shrsc_cq157;
  wire multm_reduce_mulsc_shrsc_cq158;
  wire multm_reduce_mulsc_shrsc_cq159;
  wire multm_reduce_mulsc_shrsc_cq160;
  wire multm_reduce_mulsc_shrsc_cq161;
  wire multm_reduce_mulsc_shrsc_cq162;
  wire multm_reduce_mulsc_shrsc_cq163;
  wire multm_reduce_mulsc_shrsc_cq164;
  wire multm_reduce_mulsc_shrsc_cq165;
  wire multm_reduce_mulsc_shrsc_cq166;
  wire multm_reduce_mulsc_shrsc_cq167;
  wire multm_reduce_mulsc_shrsc_cq168;
  wire multm_reduce_mulsc_shrsc_cq169;
  wire multm_reduce_mulsc_shrsc_cq170;
  wire multm_reduce_mulsc_shrsc_cq171;
  wire multm_reduce_mulsc_shrsc_cq172;
  wire multm_reduce_mulsc_shrsc_cq173;
  wire multm_reduce_mulsc_shrsc_cq174;
  wire multm_reduce_mulsc_shrsc_cq175;
  wire multm_reduce_mulsc_shrsc_cq176;
  wire multm_reduce_mulsc_shrsc_cq177;
  wire multm_reduce_mulsc_shrsc_cq178;
  wire multm_reduce_mulsc_shrsc_cq179;
  wire multm_reduce_mulsc_shrsc_cq180;
  wire multm_reduce_mulsc_shrsc_cq181;
  wire multm_reduce_mulsc_shrsc_cq182;
  wire multm_reduce_mulsc_shrsc_cr0;
  wire multm_reduce_mulsc_shrsc_cr1;
  wire multm_reduce_mulsc_shrsc_cr2;
  wire multm_reduce_mulsc_shrsc_cr3;
  wire multm_reduce_mulsc_shrsc_cr4;
  wire multm_reduce_mulsc_shrsc_cr5;
  wire multm_reduce_mulsc_shrsc_cr6;
  wire multm_reduce_mulsc_shrsc_cr7;
  wire multm_reduce_mulsc_shrsc_cr8;
  wire multm_reduce_mulsc_shrsc_cr9;
  wire multm_reduce_mulsc_shrsc_cr10;
  wire multm_reduce_mulsc_shrsc_cr11;
  wire multm_reduce_mulsc_shrsc_cr12;
  wire multm_reduce_mulsc_shrsc_cr13;
  wire multm_reduce_mulsc_shrsc_cr14;
  wire multm_reduce_mulsc_shrsc_cr15;
  wire multm_reduce_mulsc_shrsc_cr16;
  wire multm_reduce_mulsc_shrsc_cr17;
  wire multm_reduce_mulsc_shrsc_cr18;
  wire multm_reduce_mulsc_shrsc_cr19;
  wire multm_reduce_mulsc_shrsc_cr20;
  wire multm_reduce_mulsc_shrsc_cr21;
  wire multm_reduce_mulsc_shrsc_cr22;
  wire multm_reduce_mulsc_shrsc_cr23;
  wire multm_reduce_mulsc_shrsc_cr24;
  wire multm_reduce_mulsc_shrsc_cr25;
  wire multm_reduce_mulsc_shrsc_cr26;
  wire multm_reduce_mulsc_shrsc_cr27;
  wire multm_reduce_mulsc_shrsc_cr28;
  wire multm_reduce_mulsc_shrsc_cr29;
  wire multm_reduce_mulsc_shrsc_cr30;
  wire multm_reduce_mulsc_shrsc_cr31;
  wire multm_reduce_mulsc_shrsc_cr32;
  wire multm_reduce_mulsc_shrsc_cr33;
  wire multm_reduce_mulsc_shrsc_cr34;
  wire multm_reduce_mulsc_shrsc_cr35;
  wire multm_reduce_mulsc_shrsc_cr36;
  wire multm_reduce_mulsc_shrsc_cr37;
  wire multm_reduce_mulsc_shrsc_cr38;
  wire multm_reduce_mulsc_shrsc_cr39;
  wire multm_reduce_mulsc_shrsc_cr40;
  wire multm_reduce_mulsc_shrsc_cr41;
  wire multm_reduce_mulsc_shrsc_cr42;
  wire multm_reduce_mulsc_shrsc_cr43;
  wire multm_reduce_mulsc_shrsc_cr44;
  wire multm_reduce_mulsc_shrsc_cr45;
  wire multm_reduce_mulsc_shrsc_cr46;
  wire multm_reduce_mulsc_shrsc_cr47;
  wire multm_reduce_mulsc_shrsc_cr48;
  wire multm_reduce_mulsc_shrsc_cr49;
  wire multm_reduce_mulsc_shrsc_cr50;
  wire multm_reduce_mulsc_shrsc_cr51;
  wire multm_reduce_mulsc_shrsc_cr52;
  wire multm_reduce_mulsc_shrsc_cr53;
  wire multm_reduce_mulsc_shrsc_cr54;
  wire multm_reduce_mulsc_shrsc_cr55;
  wire multm_reduce_mulsc_shrsc_cr56;
  wire multm_reduce_mulsc_shrsc_cr57;
  wire multm_reduce_mulsc_shrsc_cr58;
  wire multm_reduce_mulsc_shrsc_cr59;
  wire multm_reduce_mulsc_shrsc_cr60;
  wire multm_reduce_mulsc_shrsc_cr61;
  wire multm_reduce_mulsc_shrsc_cr62;
  wire multm_reduce_mulsc_shrsc_cr63;
  wire multm_reduce_mulsc_shrsc_cr64;
  wire multm_reduce_mulsc_shrsc_cr65;
  wire multm_reduce_mulsc_shrsc_cr66;
  wire multm_reduce_mulsc_shrsc_cr67;
  wire multm_reduce_mulsc_shrsc_cr68;
  wire multm_reduce_mulsc_shrsc_cr69;
  wire multm_reduce_mulsc_shrsc_cr70;
  wire multm_reduce_mulsc_shrsc_cr71;
  wire multm_reduce_mulsc_shrsc_cr72;
  wire multm_reduce_mulsc_shrsc_cr73;
  wire multm_reduce_mulsc_shrsc_cr74;
  wire multm_reduce_mulsc_shrsc_cr75;
  wire multm_reduce_mulsc_shrsc_cr76;
  wire multm_reduce_mulsc_shrsc_cr77;
  wire multm_reduce_mulsc_shrsc_cr78;
  wire multm_reduce_mulsc_shrsc_cr79;
  wire multm_reduce_mulsc_shrsc_cr80;
  wire multm_reduce_mulsc_shrsc_cr81;
  wire multm_reduce_mulsc_shrsc_cr82;
  wire multm_reduce_mulsc_shrsc_cr83;
  wire multm_reduce_mulsc_shrsc_cr84;
  wire multm_reduce_mulsc_shrsc_cr85;
  wire multm_reduce_mulsc_shrsc_cr86;
  wire multm_reduce_mulsc_shrsc_cr87;
  wire multm_reduce_mulsc_shrsc_cr88;
  wire multm_reduce_mulsc_shrsc_cr89;
  wire multm_reduce_mulsc_shrsc_cr90;
  wire multm_reduce_mulsc_shrsc_cr91;
  wire multm_reduce_mulsc_shrsc_cr92;
  wire multm_reduce_mulsc_shrsc_cr93;
  wire multm_reduce_mulsc_shrsc_cr94;
  wire multm_reduce_mulsc_shrsc_cr95;
  wire multm_reduce_mulsc_shrsc_cr96;
  wire multm_reduce_mulsc_shrsc_cr97;
  wire multm_reduce_mulsc_shrsc_cr98;
  wire multm_reduce_mulsc_shrsc_cr99;
  wire multm_reduce_mulsc_shrsc_cr100;
  wire multm_reduce_mulsc_shrsc_cr101;
  wire multm_reduce_mulsc_shrsc_cr102;
  wire multm_reduce_mulsc_shrsc_cr103;
  wire multm_reduce_mulsc_shrsc_cr104;
  wire multm_reduce_mulsc_shrsc_cr105;
  wire multm_reduce_mulsc_shrsc_cr106;
  wire multm_reduce_mulsc_shrsc_cr107;
  wire multm_reduce_mulsc_shrsc_cr108;
  wire multm_reduce_mulsc_shrsc_cr109;
  wire multm_reduce_mulsc_shrsc_cr110;
  wire multm_reduce_mulsc_shrsc_cr111;
  wire multm_reduce_mulsc_shrsc_cr112;
  wire multm_reduce_mulsc_shrsc_cr113;
  wire multm_reduce_mulsc_shrsc_cr114;
  wire multm_reduce_mulsc_shrsc_cr115;
  wire multm_reduce_mulsc_shrsc_cr116;
  wire multm_reduce_mulsc_shrsc_cr117;
  wire multm_reduce_mulsc_shrsc_cr118;
  wire multm_reduce_mulsc_shrsc_cr119;
  wire multm_reduce_mulsc_shrsc_cr120;
  wire multm_reduce_mulsc_shrsc_cr121;
  wire multm_reduce_mulsc_shrsc_cr122;
  wire multm_reduce_mulsc_shrsc_cr123;
  wire multm_reduce_mulsc_shrsc_cr124;
  wire multm_reduce_mulsc_shrsc_cr125;
  wire multm_reduce_mulsc_shrsc_cr126;
  wire multm_reduce_mulsc_shrsc_cr127;
  wire multm_reduce_mulsc_shrsc_cr128;
  wire multm_reduce_mulsc_shrsc_cr129;
  wire multm_reduce_mulsc_shrsc_cr130;
  wire multm_reduce_mulsc_shrsc_cr131;
  wire multm_reduce_mulsc_shrsc_cr132;
  wire multm_reduce_mulsc_shrsc_cr133;
  wire multm_reduce_mulsc_shrsc_cr134;
  wire multm_reduce_mulsc_shrsc_cr135;
  wire multm_reduce_mulsc_shrsc_cr136;
  wire multm_reduce_mulsc_shrsc_cr137;
  wire multm_reduce_mulsc_shrsc_cr138;
  wire multm_reduce_mulsc_shrsc_cr139;
  wire multm_reduce_mulsc_shrsc_cr140;
  wire multm_reduce_mulsc_shrsc_cr141;
  wire multm_reduce_mulsc_shrsc_cr142;
  wire multm_reduce_mulsc_shrsc_cr143;
  wire multm_reduce_mulsc_shrsc_cr144;
  wire multm_reduce_mulsc_shrsc_cr145;
  wire multm_reduce_mulsc_shrsc_cr146;
  wire multm_reduce_mulsc_shrsc_cr147;
  wire multm_reduce_mulsc_shrsc_cr148;
  wire multm_reduce_mulsc_shrsc_cr149;
  wire multm_reduce_mulsc_shrsc_cr150;
  wire multm_reduce_mulsc_shrsc_cr151;
  wire multm_reduce_mulsc_shrsc_cr152;
  wire multm_reduce_mulsc_shrsc_cr153;
  wire multm_reduce_mulsc_shrsc_cr154;
  wire multm_reduce_mulsc_shrsc_cr155;
  wire multm_reduce_mulsc_shrsc_cr156;
  wire multm_reduce_mulsc_shrsc_cr157;
  wire multm_reduce_mulsc_shrsc_cr158;
  wire multm_reduce_mulsc_shrsc_cr159;
  wire multm_reduce_mulsc_shrsc_cr160;
  wire multm_reduce_mulsc_shrsc_cr161;
  wire multm_reduce_mulsc_shrsc_cr162;
  wire multm_reduce_mulsc_shrsc_cr163;
  wire multm_reduce_mulsc_shrsc_cr164;
  wire multm_reduce_mulsc_shrsc_cr165;
  wire multm_reduce_mulsc_shrsc_cr166;
  wire multm_reduce_mulsc_shrsc_cr167;
  wire multm_reduce_mulsc_shrsc_cr168;
  wire multm_reduce_mulsc_shrsc_cr169;
  wire multm_reduce_mulsc_shrsc_cr170;
  wire multm_reduce_mulsc_shrsc_cr171;
  wire multm_reduce_mulsc_shrsc_cr172;
  wire multm_reduce_mulsc_shrsc_cr173;
  wire multm_reduce_mulsc_shrsc_cr174;
  wire multm_reduce_mulsc_shrsc_cr175;
  wire multm_reduce_mulsc_shrsc_cr176;
  wire multm_reduce_mulsc_shrsc_cr177;
  wire multm_reduce_mulsc_shrsc_cr178;
  wire multm_reduce_mulsc_shrsc_cr179;
  wire multm_reduce_mulsc_shrsc_cr180;
  wire multm_reduce_mulsc_shrsc_cr181;
  wire multm_reduce_mulsc_shrsc_cr182;
  wire multm_reduce_mulsc_shrsc_cr183;
  wire multm_reduce_mulsc_shrsc_sq0;
  wire multm_reduce_mulsc_shrsc_sq1;
  wire multm_reduce_mulsc_shrsc_sq2;
  wire multm_reduce_mulsc_shrsc_sq3;
  wire multm_reduce_mulsc_shrsc_sq4;
  wire multm_reduce_mulsc_shrsc_sq5;
  wire multm_reduce_mulsc_shrsc_sq6;
  wire multm_reduce_mulsc_shrsc_sq7;
  wire multm_reduce_mulsc_shrsc_sq8;
  wire multm_reduce_mulsc_shrsc_sq9;
  wire multm_reduce_mulsc_shrsc_sq10;
  wire multm_reduce_mulsc_shrsc_sq11;
  wire multm_reduce_mulsc_shrsc_sq12;
  wire multm_reduce_mulsc_shrsc_sq13;
  wire multm_reduce_mulsc_shrsc_sq14;
  wire multm_reduce_mulsc_shrsc_sq15;
  wire multm_reduce_mulsc_shrsc_sq16;
  wire multm_reduce_mulsc_shrsc_sq17;
  wire multm_reduce_mulsc_shrsc_sq18;
  wire multm_reduce_mulsc_shrsc_sq19;
  wire multm_reduce_mulsc_shrsc_sq20;
  wire multm_reduce_mulsc_shrsc_sq21;
  wire multm_reduce_mulsc_shrsc_sq22;
  wire multm_reduce_mulsc_shrsc_sq23;
  wire multm_reduce_mulsc_shrsc_sq24;
  wire multm_reduce_mulsc_shrsc_sq25;
  wire multm_reduce_mulsc_shrsc_sq26;
  wire multm_reduce_mulsc_shrsc_sq27;
  wire multm_reduce_mulsc_shrsc_sq28;
  wire multm_reduce_mulsc_shrsc_sq29;
  wire multm_reduce_mulsc_shrsc_sq30;
  wire multm_reduce_mulsc_shrsc_sq31;
  wire multm_reduce_mulsc_shrsc_sq32;
  wire multm_reduce_mulsc_shrsc_sq33;
  wire multm_reduce_mulsc_shrsc_sq34;
  wire multm_reduce_mulsc_shrsc_sq35;
  wire multm_reduce_mulsc_shrsc_sq36;
  wire multm_reduce_mulsc_shrsc_sq37;
  wire multm_reduce_mulsc_shrsc_sq38;
  wire multm_reduce_mulsc_shrsc_sq39;
  wire multm_reduce_mulsc_shrsc_sq40;
  wire multm_reduce_mulsc_shrsc_sq41;
  wire multm_reduce_mulsc_shrsc_sq42;
  wire multm_reduce_mulsc_shrsc_sq43;
  wire multm_reduce_mulsc_shrsc_sq44;
  wire multm_reduce_mulsc_shrsc_sq45;
  wire multm_reduce_mulsc_shrsc_sq46;
  wire multm_reduce_mulsc_shrsc_sq47;
  wire multm_reduce_mulsc_shrsc_sq48;
  wire multm_reduce_mulsc_shrsc_sq49;
  wire multm_reduce_mulsc_shrsc_sq50;
  wire multm_reduce_mulsc_shrsc_sq51;
  wire multm_reduce_mulsc_shrsc_sq52;
  wire multm_reduce_mulsc_shrsc_sq53;
  wire multm_reduce_mulsc_shrsc_sq54;
  wire multm_reduce_mulsc_shrsc_sq55;
  wire multm_reduce_mulsc_shrsc_sq56;
  wire multm_reduce_mulsc_shrsc_sq57;
  wire multm_reduce_mulsc_shrsc_sq58;
  wire multm_reduce_mulsc_shrsc_sq59;
  wire multm_reduce_mulsc_shrsc_sq60;
  wire multm_reduce_mulsc_shrsc_sq61;
  wire multm_reduce_mulsc_shrsc_sq62;
  wire multm_reduce_mulsc_shrsc_sq63;
  wire multm_reduce_mulsc_shrsc_sq64;
  wire multm_reduce_mulsc_shrsc_sq65;
  wire multm_reduce_mulsc_shrsc_sq66;
  wire multm_reduce_mulsc_shrsc_sq67;
  wire multm_reduce_mulsc_shrsc_sq68;
  wire multm_reduce_mulsc_shrsc_sq69;
  wire multm_reduce_mulsc_shrsc_sq70;
  wire multm_reduce_mulsc_shrsc_sq71;
  wire multm_reduce_mulsc_shrsc_sq72;
  wire multm_reduce_mulsc_shrsc_sq73;
  wire multm_reduce_mulsc_shrsc_sq74;
  wire multm_reduce_mulsc_shrsc_sq75;
  wire multm_reduce_mulsc_shrsc_sq76;
  wire multm_reduce_mulsc_shrsc_sq77;
  wire multm_reduce_mulsc_shrsc_sq78;
  wire multm_reduce_mulsc_shrsc_sq79;
  wire multm_reduce_mulsc_shrsc_sq80;
  wire multm_reduce_mulsc_shrsc_sq81;
  wire multm_reduce_mulsc_shrsc_sq82;
  wire multm_reduce_mulsc_shrsc_sq83;
  wire multm_reduce_mulsc_shrsc_sq84;
  wire multm_reduce_mulsc_shrsc_sq85;
  wire multm_reduce_mulsc_shrsc_sq86;
  wire multm_reduce_mulsc_shrsc_sq87;
  wire multm_reduce_mulsc_shrsc_sq88;
  wire multm_reduce_mulsc_shrsc_sq89;
  wire multm_reduce_mulsc_shrsc_sq90;
  wire multm_reduce_mulsc_shrsc_sq91;
  wire multm_reduce_mulsc_shrsc_sq92;
  wire multm_reduce_mulsc_shrsc_sq93;
  wire multm_reduce_mulsc_shrsc_sq94;
  wire multm_reduce_mulsc_shrsc_sq95;
  wire multm_reduce_mulsc_shrsc_sq96;
  wire multm_reduce_mulsc_shrsc_sq97;
  wire multm_reduce_mulsc_shrsc_sq98;
  wire multm_reduce_mulsc_shrsc_sq99;
  wire multm_reduce_mulsc_shrsc_sq100;
  wire multm_reduce_mulsc_shrsc_sq101;
  wire multm_reduce_mulsc_shrsc_sq102;
  wire multm_reduce_mulsc_shrsc_sq103;
  wire multm_reduce_mulsc_shrsc_sq104;
  wire multm_reduce_mulsc_shrsc_sq105;
  wire multm_reduce_mulsc_shrsc_sq106;
  wire multm_reduce_mulsc_shrsc_sq107;
  wire multm_reduce_mulsc_shrsc_sq108;
  wire multm_reduce_mulsc_shrsc_sq109;
  wire multm_reduce_mulsc_shrsc_sq110;
  wire multm_reduce_mulsc_shrsc_sq111;
  wire multm_reduce_mulsc_shrsc_sq112;
  wire multm_reduce_mulsc_shrsc_sq113;
  wire multm_reduce_mulsc_shrsc_sq114;
  wire multm_reduce_mulsc_shrsc_sq115;
  wire multm_reduce_mulsc_shrsc_sq116;
  wire multm_reduce_mulsc_shrsc_sq117;
  wire multm_reduce_mulsc_shrsc_sq118;
  wire multm_reduce_mulsc_shrsc_sq119;
  wire multm_reduce_mulsc_shrsc_sq120;
  wire multm_reduce_mulsc_shrsc_sq121;
  wire multm_reduce_mulsc_shrsc_sq122;
  wire multm_reduce_mulsc_shrsc_sq123;
  wire multm_reduce_mulsc_shrsc_sq124;
  wire multm_reduce_mulsc_shrsc_sq125;
  wire multm_reduce_mulsc_shrsc_sq126;
  wire multm_reduce_mulsc_shrsc_sq127;
  wire multm_reduce_mulsc_shrsc_sq128;
  wire multm_reduce_mulsc_shrsc_sq129;
  wire multm_reduce_mulsc_shrsc_sq130;
  wire multm_reduce_mulsc_shrsc_sq131;
  wire multm_reduce_mulsc_shrsc_sq132;
  wire multm_reduce_mulsc_shrsc_sq133;
  wire multm_reduce_mulsc_shrsc_sq134;
  wire multm_reduce_mulsc_shrsc_sq135;
  wire multm_reduce_mulsc_shrsc_sq136;
  wire multm_reduce_mulsc_shrsc_sq137;
  wire multm_reduce_mulsc_shrsc_sq138;
  wire multm_reduce_mulsc_shrsc_sq139;
  wire multm_reduce_mulsc_shrsc_sq140;
  wire multm_reduce_mulsc_shrsc_sq141;
  wire multm_reduce_mulsc_shrsc_sq142;
  wire multm_reduce_mulsc_shrsc_sq143;
  wire multm_reduce_mulsc_shrsc_sq144;
  wire multm_reduce_mulsc_shrsc_sq145;
  wire multm_reduce_mulsc_shrsc_sq146;
  wire multm_reduce_mulsc_shrsc_sq147;
  wire multm_reduce_mulsc_shrsc_sq148;
  wire multm_reduce_mulsc_shrsc_sq149;
  wire multm_reduce_mulsc_shrsc_sq150;
  wire multm_reduce_mulsc_shrsc_sq151;
  wire multm_reduce_mulsc_shrsc_sq152;
  wire multm_reduce_mulsc_shrsc_sq153;
  wire multm_reduce_mulsc_shrsc_sq154;
  wire multm_reduce_mulsc_shrsc_sq155;
  wire multm_reduce_mulsc_shrsc_sq156;
  wire multm_reduce_mulsc_shrsc_sq157;
  wire multm_reduce_mulsc_shrsc_sq158;
  wire multm_reduce_mulsc_shrsc_sq159;
  wire multm_reduce_mulsc_shrsc_sq160;
  wire multm_reduce_mulsc_shrsc_sq161;
  wire multm_reduce_mulsc_shrsc_sq162;
  wire multm_reduce_mulsc_shrsc_sq163;
  wire multm_reduce_mulsc_shrsc_sq164;
  wire multm_reduce_mulsc_shrsc_sq165;
  wire multm_reduce_mulsc_shrsc_sq166;
  wire multm_reduce_mulsc_shrsc_sq167;
  wire multm_reduce_mulsc_shrsc_sq168;
  wire multm_reduce_mulsc_shrsc_sq169;
  wire multm_reduce_mulsc_shrsc_sq170;
  wire multm_reduce_mulsc_shrsc_sq171;
  wire multm_reduce_mulsc_shrsc_sq172;
  wire multm_reduce_mulsc_shrsc_sq173;
  wire multm_reduce_mulsc_shrsc_sq174;
  wire multm_reduce_mulsc_shrsc_sq175;
  wire multm_reduce_mulsc_shrsc_sq176;
  wire multm_reduce_mulsc_shrsc_sq177;
  wire multm_reduce_mulsc_shrsc_sq178;
  wire multm_reduce_mulsc_shrsc_sq179;
  wire multm_reduce_mulsc_shrsc_sq180;
  wire multm_reduce_mulsc_shrsc_sq181;
  wire multm_reduce_mulsc_shrsc_sq182;
  wire multm_reduce_mulsc_shrsc_sr0;
  wire multm_reduce_mulsc_shrsc_sr1;
  wire multm_reduce_mulsc_shrsc_sr2;
  wire multm_reduce_mulsc_shrsc_sr3;
  wire multm_reduce_mulsc_shrsc_sr4;
  wire multm_reduce_mulsc_shrsc_sr5;
  wire multm_reduce_mulsc_shrsc_sr6;
  wire multm_reduce_mulsc_shrsc_sr7;
  wire multm_reduce_mulsc_shrsc_sr8;
  wire multm_reduce_mulsc_shrsc_sr9;
  wire multm_reduce_mulsc_shrsc_sr10;
  wire multm_reduce_mulsc_shrsc_sr11;
  wire multm_reduce_mulsc_shrsc_sr12;
  wire multm_reduce_mulsc_shrsc_sr13;
  wire multm_reduce_mulsc_shrsc_sr14;
  wire multm_reduce_mulsc_shrsc_sr15;
  wire multm_reduce_mulsc_shrsc_sr16;
  wire multm_reduce_mulsc_shrsc_sr17;
  wire multm_reduce_mulsc_shrsc_sr18;
  wire multm_reduce_mulsc_shrsc_sr19;
  wire multm_reduce_mulsc_shrsc_sr20;
  wire multm_reduce_mulsc_shrsc_sr21;
  wire multm_reduce_mulsc_shrsc_sr22;
  wire multm_reduce_mulsc_shrsc_sr23;
  wire multm_reduce_mulsc_shrsc_sr24;
  wire multm_reduce_mulsc_shrsc_sr25;
  wire multm_reduce_mulsc_shrsc_sr26;
  wire multm_reduce_mulsc_shrsc_sr27;
  wire multm_reduce_mulsc_shrsc_sr28;
  wire multm_reduce_mulsc_shrsc_sr29;
  wire multm_reduce_mulsc_shrsc_sr30;
  wire multm_reduce_mulsc_shrsc_sr31;
  wire multm_reduce_mulsc_shrsc_sr32;
  wire multm_reduce_mulsc_shrsc_sr33;
  wire multm_reduce_mulsc_shrsc_sr34;
  wire multm_reduce_mulsc_shrsc_sr35;
  wire multm_reduce_mulsc_shrsc_sr36;
  wire multm_reduce_mulsc_shrsc_sr37;
  wire multm_reduce_mulsc_shrsc_sr38;
  wire multm_reduce_mulsc_shrsc_sr39;
  wire multm_reduce_mulsc_shrsc_sr40;
  wire multm_reduce_mulsc_shrsc_sr41;
  wire multm_reduce_mulsc_shrsc_sr42;
  wire multm_reduce_mulsc_shrsc_sr43;
  wire multm_reduce_mulsc_shrsc_sr44;
  wire multm_reduce_mulsc_shrsc_sr45;
  wire multm_reduce_mulsc_shrsc_sr46;
  wire multm_reduce_mulsc_shrsc_sr47;
  wire multm_reduce_mulsc_shrsc_sr48;
  wire multm_reduce_mulsc_shrsc_sr49;
  wire multm_reduce_mulsc_shrsc_sr50;
  wire multm_reduce_mulsc_shrsc_sr51;
  wire multm_reduce_mulsc_shrsc_sr52;
  wire multm_reduce_mulsc_shrsc_sr53;
  wire multm_reduce_mulsc_shrsc_sr54;
  wire multm_reduce_mulsc_shrsc_sr55;
  wire multm_reduce_mulsc_shrsc_sr56;
  wire multm_reduce_mulsc_shrsc_sr57;
  wire multm_reduce_mulsc_shrsc_sr58;
  wire multm_reduce_mulsc_shrsc_sr59;
  wire multm_reduce_mulsc_shrsc_sr60;
  wire multm_reduce_mulsc_shrsc_sr61;
  wire multm_reduce_mulsc_shrsc_sr62;
  wire multm_reduce_mulsc_shrsc_sr63;
  wire multm_reduce_mulsc_shrsc_sr64;
  wire multm_reduce_mulsc_shrsc_sr65;
  wire multm_reduce_mulsc_shrsc_sr66;
  wire multm_reduce_mulsc_shrsc_sr67;
  wire multm_reduce_mulsc_shrsc_sr68;
  wire multm_reduce_mulsc_shrsc_sr69;
  wire multm_reduce_mulsc_shrsc_sr70;
  wire multm_reduce_mulsc_shrsc_sr71;
  wire multm_reduce_mulsc_shrsc_sr72;
  wire multm_reduce_mulsc_shrsc_sr73;
  wire multm_reduce_mulsc_shrsc_sr74;
  wire multm_reduce_mulsc_shrsc_sr75;
  wire multm_reduce_mulsc_shrsc_sr76;
  wire multm_reduce_mulsc_shrsc_sr77;
  wire multm_reduce_mulsc_shrsc_sr78;
  wire multm_reduce_mulsc_shrsc_sr79;
  wire multm_reduce_mulsc_shrsc_sr80;
  wire multm_reduce_mulsc_shrsc_sr81;
  wire multm_reduce_mulsc_shrsc_sr82;
  wire multm_reduce_mulsc_shrsc_sr83;
  wire multm_reduce_mulsc_shrsc_sr84;
  wire multm_reduce_mulsc_shrsc_sr85;
  wire multm_reduce_mulsc_shrsc_sr86;
  wire multm_reduce_mulsc_shrsc_sr87;
  wire multm_reduce_mulsc_shrsc_sr88;
  wire multm_reduce_mulsc_shrsc_sr89;
  wire multm_reduce_mulsc_shrsc_sr90;
  wire multm_reduce_mulsc_shrsc_sr91;
  wire multm_reduce_mulsc_shrsc_sr92;
  wire multm_reduce_mulsc_shrsc_sr93;
  wire multm_reduce_mulsc_shrsc_sr94;
  wire multm_reduce_mulsc_shrsc_sr95;
  wire multm_reduce_mulsc_shrsc_sr96;
  wire multm_reduce_mulsc_shrsc_sr97;
  wire multm_reduce_mulsc_shrsc_sr98;
  wire multm_reduce_mulsc_shrsc_sr99;
  wire multm_reduce_mulsc_shrsc_sr100;
  wire multm_reduce_mulsc_shrsc_sr101;
  wire multm_reduce_mulsc_shrsc_sr102;
  wire multm_reduce_mulsc_shrsc_sr103;
  wire multm_reduce_mulsc_shrsc_sr104;
  wire multm_reduce_mulsc_shrsc_sr105;
  wire multm_reduce_mulsc_shrsc_sr106;
  wire multm_reduce_mulsc_shrsc_sr107;
  wire multm_reduce_mulsc_shrsc_sr108;
  wire multm_reduce_mulsc_shrsc_sr109;
  wire multm_reduce_mulsc_shrsc_sr110;
  wire multm_reduce_mulsc_shrsc_sr111;
  wire multm_reduce_mulsc_shrsc_sr112;
  wire multm_reduce_mulsc_shrsc_sr113;
  wire multm_reduce_mulsc_shrsc_sr114;
  wire multm_reduce_mulsc_shrsc_sr115;
  wire multm_reduce_mulsc_shrsc_sr116;
  wire multm_reduce_mulsc_shrsc_sr117;
  wire multm_reduce_mulsc_shrsc_sr118;
  wire multm_reduce_mulsc_shrsc_sr119;
  wire multm_reduce_mulsc_shrsc_sr120;
  wire multm_reduce_mulsc_shrsc_sr121;
  wire multm_reduce_mulsc_shrsc_sr122;
  wire multm_reduce_mulsc_shrsc_sr123;
  wire multm_reduce_mulsc_shrsc_sr124;
  wire multm_reduce_mulsc_shrsc_sr125;
  wire multm_reduce_mulsc_shrsc_sr126;
  wire multm_reduce_mulsc_shrsc_sr127;
  wire multm_reduce_mulsc_shrsc_sr128;
  wire multm_reduce_mulsc_shrsc_sr129;
  wire multm_reduce_mulsc_shrsc_sr130;
  wire multm_reduce_mulsc_shrsc_sr131;
  wire multm_reduce_mulsc_shrsc_sr132;
  wire multm_reduce_mulsc_shrsc_sr133;
  wire multm_reduce_mulsc_shrsc_sr134;
  wire multm_reduce_mulsc_shrsc_sr135;
  wire multm_reduce_mulsc_shrsc_sr136;
  wire multm_reduce_mulsc_shrsc_sr137;
  wire multm_reduce_mulsc_shrsc_sr138;
  wire multm_reduce_mulsc_shrsc_sr139;
  wire multm_reduce_mulsc_shrsc_sr140;
  wire multm_reduce_mulsc_shrsc_sr141;
  wire multm_reduce_mulsc_shrsc_sr142;
  wire multm_reduce_mulsc_shrsc_sr143;
  wire multm_reduce_mulsc_shrsc_sr144;
  wire multm_reduce_mulsc_shrsc_sr145;
  wire multm_reduce_mulsc_shrsc_sr146;
  wire multm_reduce_mulsc_shrsc_sr147;
  wire multm_reduce_mulsc_shrsc_sr148;
  wire multm_reduce_mulsc_shrsc_sr149;
  wire multm_reduce_mulsc_shrsc_sr150;
  wire multm_reduce_mulsc_shrsc_sr151;
  wire multm_reduce_mulsc_shrsc_sr152;
  wire multm_reduce_mulsc_shrsc_sr153;
  wire multm_reduce_mulsc_shrsc_sr154;
  wire multm_reduce_mulsc_shrsc_sr155;
  wire multm_reduce_mulsc_shrsc_sr156;
  wire multm_reduce_mulsc_shrsc_sr157;
  wire multm_reduce_mulsc_shrsc_sr158;
  wire multm_reduce_mulsc_shrsc_sr159;
  wire multm_reduce_mulsc_shrsc_sr160;
  wire multm_reduce_mulsc_shrsc_sr161;
  wire multm_reduce_mulsc_shrsc_sr162;
  wire multm_reduce_mulsc_shrsc_sr163;
  wire multm_reduce_mulsc_shrsc_sr164;
  wire multm_reduce_mulsc_shrsc_sr165;
  wire multm_reduce_mulsc_shrsc_sr166;
  wire multm_reduce_mulsc_shrsc_sr167;
  wire multm_reduce_mulsc_shrsc_sr168;
  wire multm_reduce_mulsc_shrsc_sr169;
  wire multm_reduce_mulsc_shrsc_sr170;
  wire multm_reduce_mulsc_shrsc_sr171;
  wire multm_reduce_mulsc_shrsc_sr172;
  wire multm_reduce_mulsc_shrsc_sr173;
  wire multm_reduce_mulsc_shrsc_sr174;
  wire multm_reduce_mulsc_shrsc_sr175;
  wire multm_reduce_mulsc_shrsc_sr176;
  wire multm_reduce_mulsc_shrsc_sr177;
  wire multm_reduce_mulsc_shrsc_sr178;
  wire multm_reduce_mulsc_shrsc_sr179;
  wire multm_reduce_mulsc_shrsc_sr180;
  wire multm_reduce_mulsc_shrsc_sr181;
  wire multm_reduce_mulsc_shrsc_sr182;
  wire multm_reduce_mulsc_xb;
  wire multm_reduce_mw;
  wire multm_reduce_or3_wx;
  wire multm_reduce_pb;
  wire multm_reduce_pc0;
  wire multm_reduce_pc1;
  wire multm_reduce_pc2;
  wire multm_reduce_pc3;
  wire multm_reduce_pc4;
  wire multm_reduce_pc5;
  wire multm_reduce_pc6;
  wire multm_reduce_pc7;
  wire multm_reduce_pc8;
  wire multm_reduce_pc9;
  wire multm_reduce_pc10;
  wire multm_reduce_pc11;
  wire multm_reduce_pc12;
  wire multm_reduce_pc13;
  wire multm_reduce_pc14;
  wire multm_reduce_pc15;
  wire multm_reduce_pc16;
  wire multm_reduce_pc17;
  wire multm_reduce_pc18;
  wire multm_reduce_pc19;
  wire multm_reduce_pc20;
  wire multm_reduce_pc21;
  wire multm_reduce_pc22;
  wire multm_reduce_pc23;
  wire multm_reduce_pc24;
  wire multm_reduce_pc25;
  wire multm_reduce_pc26;
  wire multm_reduce_pc27;
  wire multm_reduce_pc28;
  wire multm_reduce_pc29;
  wire multm_reduce_pc30;
  wire multm_reduce_pc31;
  wire multm_reduce_pc32;
  wire multm_reduce_pc33;
  wire multm_reduce_pc34;
  wire multm_reduce_pc35;
  wire multm_reduce_pc36;
  wire multm_reduce_pc37;
  wire multm_reduce_pc38;
  wire multm_reduce_pc39;
  wire multm_reduce_pc40;
  wire multm_reduce_pc41;
  wire multm_reduce_pc42;
  wire multm_reduce_pc43;
  wire multm_reduce_pc44;
  wire multm_reduce_pc45;
  wire multm_reduce_pc46;
  wire multm_reduce_pc47;
  wire multm_reduce_pc48;
  wire multm_reduce_pc49;
  wire multm_reduce_pc50;
  wire multm_reduce_pc51;
  wire multm_reduce_pc52;
  wire multm_reduce_pc53;
  wire multm_reduce_pc54;
  wire multm_reduce_pc55;
  wire multm_reduce_pc56;
  wire multm_reduce_pc57;
  wire multm_reduce_pc58;
  wire multm_reduce_pc59;
  wire multm_reduce_pc60;
  wire multm_reduce_pc61;
  wire multm_reduce_pc62;
  wire multm_reduce_pc63;
  wire multm_reduce_pc64;
  wire multm_reduce_pc65;
  wire multm_reduce_pc66;
  wire multm_reduce_pc67;
  wire multm_reduce_pc68;
  wire multm_reduce_pc69;
  wire multm_reduce_pc70;
  wire multm_reduce_pc71;
  wire multm_reduce_pc72;
  wire multm_reduce_pc73;
  wire multm_reduce_pc74;
  wire multm_reduce_pc75;
  wire multm_reduce_pc76;
  wire multm_reduce_pc77;
  wire multm_reduce_pc78;
  wire multm_reduce_pc79;
  wire multm_reduce_pc80;
  wire multm_reduce_pc81;
  wire multm_reduce_pc82;
  wire multm_reduce_pc83;
  wire multm_reduce_pc84;
  wire multm_reduce_pc85;
  wire multm_reduce_pc86;
  wire multm_reduce_pc87;
  wire multm_reduce_pc88;
  wire multm_reduce_pc89;
  wire multm_reduce_pc90;
  wire multm_reduce_pc91;
  wire multm_reduce_pc92;
  wire multm_reduce_pc93;
  wire multm_reduce_pc94;
  wire multm_reduce_pc95;
  wire multm_reduce_pc96;
  wire multm_reduce_pc97;
  wire multm_reduce_pc98;
  wire multm_reduce_pc99;
  wire multm_reduce_pc100;
  wire multm_reduce_pc101;
  wire multm_reduce_pc102;
  wire multm_reduce_pc103;
  wire multm_reduce_pc104;
  wire multm_reduce_pc105;
  wire multm_reduce_pc106;
  wire multm_reduce_pc107;
  wire multm_reduce_pc108;
  wire multm_reduce_pc109;
  wire multm_reduce_pc110;
  wire multm_reduce_pc111;
  wire multm_reduce_pc112;
  wire multm_reduce_pc113;
  wire multm_reduce_pc114;
  wire multm_reduce_pc115;
  wire multm_reduce_pc116;
  wire multm_reduce_pc117;
  wire multm_reduce_pc118;
  wire multm_reduce_pc119;
  wire multm_reduce_pc120;
  wire multm_reduce_pc121;
  wire multm_reduce_pc122;
  wire multm_reduce_pc123;
  wire multm_reduce_pc124;
  wire multm_reduce_pc125;
  wire multm_reduce_pc126;
  wire multm_reduce_pc127;
  wire multm_reduce_pc128;
  wire multm_reduce_pc129;
  wire multm_reduce_pc130;
  wire multm_reduce_pc131;
  wire multm_reduce_pc132;
  wire multm_reduce_pc133;
  wire multm_reduce_pc134;
  wire multm_reduce_pc135;
  wire multm_reduce_pc136;
  wire multm_reduce_pc137;
  wire multm_reduce_pc138;
  wire multm_reduce_pc139;
  wire multm_reduce_pc140;
  wire multm_reduce_pc141;
  wire multm_reduce_pc142;
  wire multm_reduce_pc143;
  wire multm_reduce_pc144;
  wire multm_reduce_pc145;
  wire multm_reduce_pc146;
  wire multm_reduce_pc147;
  wire multm_reduce_pc148;
  wire multm_reduce_pc149;
  wire multm_reduce_pc150;
  wire multm_reduce_pc151;
  wire multm_reduce_pc152;
  wire multm_reduce_pc153;
  wire multm_reduce_pc154;
  wire multm_reduce_pc155;
  wire multm_reduce_pc156;
  wire multm_reduce_pc157;
  wire multm_reduce_pc158;
  wire multm_reduce_pc159;
  wire multm_reduce_pc160;
  wire multm_reduce_pc161;
  wire multm_reduce_pc162;
  wire multm_reduce_pc163;
  wire multm_reduce_pc164;
  wire multm_reduce_pc165;
  wire multm_reduce_pc166;
  wire multm_reduce_pc167;
  wire multm_reduce_pc168;
  wire multm_reduce_pc169;
  wire multm_reduce_pc170;
  wire multm_reduce_pc171;
  wire multm_reduce_pc172;
  wire multm_reduce_pc173;
  wire multm_reduce_pc174;
  wire multm_reduce_pc175;
  wire multm_reduce_pc176;
  wire multm_reduce_pc177;
  wire multm_reduce_pc178;
  wire multm_reduce_pc179;
  wire multm_reduce_pc180;
  wire multm_reduce_pc181;
  wire multm_reduce_pc182;
  wire multm_reduce_pc183;
  wire multm_reduce_ps0;
  wire multm_reduce_ps1;
  wire multm_reduce_ps2;
  wire multm_reduce_ps3;
  wire multm_reduce_ps4;
  wire multm_reduce_ps5;
  wire multm_reduce_ps6;
  wire multm_reduce_ps7;
  wire multm_reduce_ps8;
  wire multm_reduce_ps9;
  wire multm_reduce_ps10;
  wire multm_reduce_ps11;
  wire multm_reduce_ps12;
  wire multm_reduce_ps13;
  wire multm_reduce_ps14;
  wire multm_reduce_ps15;
  wire multm_reduce_ps16;
  wire multm_reduce_ps17;
  wire multm_reduce_ps18;
  wire multm_reduce_ps19;
  wire multm_reduce_ps20;
  wire multm_reduce_ps21;
  wire multm_reduce_ps22;
  wire multm_reduce_ps23;
  wire multm_reduce_ps24;
  wire multm_reduce_ps25;
  wire multm_reduce_ps26;
  wire multm_reduce_ps27;
  wire multm_reduce_ps28;
  wire multm_reduce_ps29;
  wire multm_reduce_ps30;
  wire multm_reduce_ps31;
  wire multm_reduce_ps32;
  wire multm_reduce_ps33;
  wire multm_reduce_ps34;
  wire multm_reduce_ps35;
  wire multm_reduce_ps36;
  wire multm_reduce_ps37;
  wire multm_reduce_ps38;
  wire multm_reduce_ps39;
  wire multm_reduce_ps40;
  wire multm_reduce_ps41;
  wire multm_reduce_ps42;
  wire multm_reduce_ps43;
  wire multm_reduce_ps44;
  wire multm_reduce_ps45;
  wire multm_reduce_ps46;
  wire multm_reduce_ps47;
  wire multm_reduce_ps48;
  wire multm_reduce_ps49;
  wire multm_reduce_ps50;
  wire multm_reduce_ps51;
  wire multm_reduce_ps52;
  wire multm_reduce_ps53;
  wire multm_reduce_ps54;
  wire multm_reduce_ps55;
  wire multm_reduce_ps56;
  wire multm_reduce_ps57;
  wire multm_reduce_ps58;
  wire multm_reduce_ps59;
  wire multm_reduce_ps60;
  wire multm_reduce_ps61;
  wire multm_reduce_ps62;
  wire multm_reduce_ps63;
  wire multm_reduce_ps64;
  wire multm_reduce_ps65;
  wire multm_reduce_ps66;
  wire multm_reduce_ps67;
  wire multm_reduce_ps68;
  wire multm_reduce_ps69;
  wire multm_reduce_ps70;
  wire multm_reduce_ps71;
  wire multm_reduce_ps72;
  wire multm_reduce_ps73;
  wire multm_reduce_ps74;
  wire multm_reduce_ps75;
  wire multm_reduce_ps76;
  wire multm_reduce_ps77;
  wire multm_reduce_ps78;
  wire multm_reduce_ps79;
  wire multm_reduce_ps80;
  wire multm_reduce_ps81;
  wire multm_reduce_ps82;
  wire multm_reduce_ps83;
  wire multm_reduce_ps84;
  wire multm_reduce_ps85;
  wire multm_reduce_ps86;
  wire multm_reduce_ps87;
  wire multm_reduce_ps88;
  wire multm_reduce_ps89;
  wire multm_reduce_ps90;
  wire multm_reduce_ps91;
  wire multm_reduce_ps92;
  wire multm_reduce_ps93;
  wire multm_reduce_ps94;
  wire multm_reduce_ps95;
  wire multm_reduce_ps96;
  wire multm_reduce_ps97;
  wire multm_reduce_ps98;
  wire multm_reduce_ps99;
  wire multm_reduce_ps100;
  wire multm_reduce_ps101;
  wire multm_reduce_ps102;
  wire multm_reduce_ps103;
  wire multm_reduce_ps104;
  wire multm_reduce_ps105;
  wire multm_reduce_ps106;
  wire multm_reduce_ps107;
  wire multm_reduce_ps108;
  wire multm_reduce_ps109;
  wire multm_reduce_ps110;
  wire multm_reduce_ps111;
  wire multm_reduce_ps112;
  wire multm_reduce_ps113;
  wire multm_reduce_ps114;
  wire multm_reduce_ps115;
  wire multm_reduce_ps116;
  wire multm_reduce_ps117;
  wire multm_reduce_ps118;
  wire multm_reduce_ps119;
  wire multm_reduce_ps120;
  wire multm_reduce_ps121;
  wire multm_reduce_ps122;
  wire multm_reduce_ps123;
  wire multm_reduce_ps124;
  wire multm_reduce_ps125;
  wire multm_reduce_ps126;
  wire multm_reduce_ps127;
  wire multm_reduce_ps128;
  wire multm_reduce_ps129;
  wire multm_reduce_ps130;
  wire multm_reduce_ps131;
  wire multm_reduce_ps132;
  wire multm_reduce_ps133;
  wire multm_reduce_ps134;
  wire multm_reduce_ps135;
  wire multm_reduce_ps136;
  wire multm_reduce_ps137;
  wire multm_reduce_ps138;
  wire multm_reduce_ps139;
  wire multm_reduce_ps140;
  wire multm_reduce_ps141;
  wire multm_reduce_ps142;
  wire multm_reduce_ps143;
  wire multm_reduce_ps144;
  wire multm_reduce_ps145;
  wire multm_reduce_ps146;
  wire multm_reduce_ps147;
  wire multm_reduce_ps148;
  wire multm_reduce_ps149;
  wire multm_reduce_ps150;
  wire multm_reduce_ps151;
  wire multm_reduce_ps152;
  wire multm_reduce_ps153;
  wire multm_reduce_ps154;
  wire multm_reduce_ps155;
  wire multm_reduce_ps156;
  wire multm_reduce_ps157;
  wire multm_reduce_ps158;
  wire multm_reduce_ps159;
  wire multm_reduce_ps160;
  wire multm_reduce_ps161;
  wire multm_reduce_ps162;
  wire multm_reduce_ps163;
  wire multm_reduce_ps164;
  wire multm_reduce_ps165;
  wire multm_reduce_ps166;
  wire multm_reduce_ps167;
  wire multm_reduce_ps168;
  wire multm_reduce_ps169;
  wire multm_reduce_ps170;
  wire multm_reduce_ps171;
  wire multm_reduce_ps172;
  wire multm_reduce_ps173;
  wire multm_reduce_ps174;
  wire multm_reduce_ps175;
  wire multm_reduce_ps176;
  wire multm_reduce_ps177;
  wire multm_reduce_ps178;
  wire multm_reduce_ps179;
  wire multm_reduce_ps180;
  wire multm_reduce_ps181;
  wire multm_reduce_ps182;
  wire multm_reduce_ps183;
  wire multm_reduce_qb;
  wire multm_reduce_qc0;
  wire multm_reduce_qc1;
  wire multm_reduce_qc2;
  wire multm_reduce_qc3;
  wire multm_reduce_qc4;
  wire multm_reduce_qc5;
  wire multm_reduce_qc6;
  wire multm_reduce_qc7;
  wire multm_reduce_qc8;
  wire multm_reduce_qc9;
  wire multm_reduce_qc10;
  wire multm_reduce_qc11;
  wire multm_reduce_qc12;
  wire multm_reduce_qc13;
  wire multm_reduce_qc14;
  wire multm_reduce_qc15;
  wire multm_reduce_qc16;
  wire multm_reduce_qc17;
  wire multm_reduce_qc18;
  wire multm_reduce_qc19;
  wire multm_reduce_qc20;
  wire multm_reduce_qc21;
  wire multm_reduce_qc22;
  wire multm_reduce_qc23;
  wire multm_reduce_qc24;
  wire multm_reduce_qc25;
  wire multm_reduce_qc26;
  wire multm_reduce_qc27;
  wire multm_reduce_qc28;
  wire multm_reduce_qc29;
  wire multm_reduce_qc30;
  wire multm_reduce_qc31;
  wire multm_reduce_qc32;
  wire multm_reduce_qc33;
  wire multm_reduce_qc34;
  wire multm_reduce_qc35;
  wire multm_reduce_qc36;
  wire multm_reduce_qc37;
  wire multm_reduce_qc38;
  wire multm_reduce_qc39;
  wire multm_reduce_qc40;
  wire multm_reduce_qc41;
  wire multm_reduce_qc42;
  wire multm_reduce_qc43;
  wire multm_reduce_qc44;
  wire multm_reduce_qc45;
  wire multm_reduce_qc46;
  wire multm_reduce_qc47;
  wire multm_reduce_qc48;
  wire multm_reduce_qc49;
  wire multm_reduce_qc50;
  wire multm_reduce_qc51;
  wire multm_reduce_qc52;
  wire multm_reduce_qc53;
  wire multm_reduce_qc54;
  wire multm_reduce_qc55;
  wire multm_reduce_qc56;
  wire multm_reduce_qc57;
  wire multm_reduce_qc58;
  wire multm_reduce_qc59;
  wire multm_reduce_qc60;
  wire multm_reduce_qc61;
  wire multm_reduce_qc62;
  wire multm_reduce_qc63;
  wire multm_reduce_qc64;
  wire multm_reduce_qc65;
  wire multm_reduce_qc66;
  wire multm_reduce_qc67;
  wire multm_reduce_qc68;
  wire multm_reduce_qc69;
  wire multm_reduce_qc70;
  wire multm_reduce_qc71;
  wire multm_reduce_qc72;
  wire multm_reduce_qc73;
  wire multm_reduce_qc74;
  wire multm_reduce_qc75;
  wire multm_reduce_qc76;
  wire multm_reduce_qc77;
  wire multm_reduce_qc78;
  wire multm_reduce_qc79;
  wire multm_reduce_qc80;
  wire multm_reduce_qc81;
  wire multm_reduce_qc82;
  wire multm_reduce_qc83;
  wire multm_reduce_qc84;
  wire multm_reduce_qc85;
  wire multm_reduce_qc86;
  wire multm_reduce_qc87;
  wire multm_reduce_qc88;
  wire multm_reduce_qc89;
  wire multm_reduce_qc90;
  wire multm_reduce_qc91;
  wire multm_reduce_qc92;
  wire multm_reduce_qc93;
  wire multm_reduce_qc94;
  wire multm_reduce_qc95;
  wire multm_reduce_qc96;
  wire multm_reduce_qc97;
  wire multm_reduce_qc98;
  wire multm_reduce_qc99;
  wire multm_reduce_qc100;
  wire multm_reduce_qc101;
  wire multm_reduce_qc102;
  wire multm_reduce_qc103;
  wire multm_reduce_qc104;
  wire multm_reduce_qc105;
  wire multm_reduce_qc106;
  wire multm_reduce_qc107;
  wire multm_reduce_qc108;
  wire multm_reduce_qc109;
  wire multm_reduce_qc110;
  wire multm_reduce_qc111;
  wire multm_reduce_qc112;
  wire multm_reduce_qc113;
  wire multm_reduce_qc114;
  wire multm_reduce_qc115;
  wire multm_reduce_qc116;
  wire multm_reduce_qc117;
  wire multm_reduce_qc118;
  wire multm_reduce_qc119;
  wire multm_reduce_qc120;
  wire multm_reduce_qc121;
  wire multm_reduce_qc122;
  wire multm_reduce_qc123;
  wire multm_reduce_qc124;
  wire multm_reduce_qc125;
  wire multm_reduce_qc126;
  wire multm_reduce_qc127;
  wire multm_reduce_qc128;
  wire multm_reduce_qc129;
  wire multm_reduce_qc130;
  wire multm_reduce_qc131;
  wire multm_reduce_qc132;
  wire multm_reduce_qc133;
  wire multm_reduce_qc134;
  wire multm_reduce_qc135;
  wire multm_reduce_qc136;
  wire multm_reduce_qc137;
  wire multm_reduce_qc138;
  wire multm_reduce_qc139;
  wire multm_reduce_qc140;
  wire multm_reduce_qc141;
  wire multm_reduce_qc142;
  wire multm_reduce_qc143;
  wire multm_reduce_qc144;
  wire multm_reduce_qc145;
  wire multm_reduce_qc146;
  wire multm_reduce_qc147;
  wire multm_reduce_qc148;
  wire multm_reduce_qc149;
  wire multm_reduce_qc150;
  wire multm_reduce_qc151;
  wire multm_reduce_qc152;
  wire multm_reduce_qc153;
  wire multm_reduce_qc154;
  wire multm_reduce_qc155;
  wire multm_reduce_qc156;
  wire multm_reduce_qc157;
  wire multm_reduce_qc158;
  wire multm_reduce_qc159;
  wire multm_reduce_qc160;
  wire multm_reduce_qc161;
  wire multm_reduce_qc162;
  wire multm_reduce_qc163;
  wire multm_reduce_qc164;
  wire multm_reduce_qc165;
  wire multm_reduce_qc166;
  wire multm_reduce_qc167;
  wire multm_reduce_qc168;
  wire multm_reduce_qc169;
  wire multm_reduce_qc170;
  wire multm_reduce_qc171;
  wire multm_reduce_qc172;
  wire multm_reduce_qc173;
  wire multm_reduce_qc174;
  wire multm_reduce_qc175;
  wire multm_reduce_qc176;
  wire multm_reduce_qc177;
  wire multm_reduce_qc178;
  wire multm_reduce_qc179;
  wire multm_reduce_qc180;
  wire multm_reduce_qc181;
  wire multm_reduce_qc182;
  wire multm_reduce_qc183;
  wire multm_reduce_qc184;
  wire multm_reduce_qs0;
  wire multm_reduce_qs1;
  wire multm_reduce_qs2;
  wire multm_reduce_qs3;
  wire multm_reduce_qs4;
  wire multm_reduce_qs5;
  wire multm_reduce_qs6;
  wire multm_reduce_qs7;
  wire multm_reduce_qs8;
  wire multm_reduce_qs9;
  wire multm_reduce_qs10;
  wire multm_reduce_qs11;
  wire multm_reduce_qs12;
  wire multm_reduce_qs13;
  wire multm_reduce_qs14;
  wire multm_reduce_qs15;
  wire multm_reduce_qs16;
  wire multm_reduce_qs17;
  wire multm_reduce_qs18;
  wire multm_reduce_qs19;
  wire multm_reduce_qs20;
  wire multm_reduce_qs21;
  wire multm_reduce_qs22;
  wire multm_reduce_qs23;
  wire multm_reduce_qs24;
  wire multm_reduce_qs25;
  wire multm_reduce_qs26;
  wire multm_reduce_qs27;
  wire multm_reduce_qs28;
  wire multm_reduce_qs29;
  wire multm_reduce_qs30;
  wire multm_reduce_qs31;
  wire multm_reduce_qs32;
  wire multm_reduce_qs33;
  wire multm_reduce_qs34;
  wire multm_reduce_qs35;
  wire multm_reduce_qs36;
  wire multm_reduce_qs37;
  wire multm_reduce_qs38;
  wire multm_reduce_qs39;
  wire multm_reduce_qs40;
  wire multm_reduce_qs41;
  wire multm_reduce_qs42;
  wire multm_reduce_qs43;
  wire multm_reduce_qs44;
  wire multm_reduce_qs45;
  wire multm_reduce_qs46;
  wire multm_reduce_qs47;
  wire multm_reduce_qs48;
  wire multm_reduce_qs49;
  wire multm_reduce_qs50;
  wire multm_reduce_qs51;
  wire multm_reduce_qs52;
  wire multm_reduce_qs53;
  wire multm_reduce_qs54;
  wire multm_reduce_qs55;
  wire multm_reduce_qs56;
  wire multm_reduce_qs57;
  wire multm_reduce_qs58;
  wire multm_reduce_qs59;
  wire multm_reduce_qs60;
  wire multm_reduce_qs61;
  wire multm_reduce_qs62;
  wire multm_reduce_qs63;
  wire multm_reduce_qs64;
  wire multm_reduce_qs65;
  wire multm_reduce_qs66;
  wire multm_reduce_qs67;
  wire multm_reduce_qs68;
  wire multm_reduce_qs69;
  wire multm_reduce_qs70;
  wire multm_reduce_qs71;
  wire multm_reduce_qs72;
  wire multm_reduce_qs73;
  wire multm_reduce_qs74;
  wire multm_reduce_qs75;
  wire multm_reduce_qs76;
  wire multm_reduce_qs77;
  wire multm_reduce_qs78;
  wire multm_reduce_qs79;
  wire multm_reduce_qs80;
  wire multm_reduce_qs81;
  wire multm_reduce_qs82;
  wire multm_reduce_qs83;
  wire multm_reduce_qs84;
  wire multm_reduce_qs85;
  wire multm_reduce_qs86;
  wire multm_reduce_qs87;
  wire multm_reduce_qs88;
  wire multm_reduce_qs89;
  wire multm_reduce_qs90;
  wire multm_reduce_qs91;
  wire multm_reduce_qs92;
  wire multm_reduce_qs93;
  wire multm_reduce_qs94;
  wire multm_reduce_qs95;
  wire multm_reduce_qs96;
  wire multm_reduce_qs97;
  wire multm_reduce_qs98;
  wire multm_reduce_qs99;
  wire multm_reduce_qs100;
  wire multm_reduce_qs101;
  wire multm_reduce_qs102;
  wire multm_reduce_qs103;
  wire multm_reduce_qs104;
  wire multm_reduce_qs105;
  wire multm_reduce_qs106;
  wire multm_reduce_qs107;
  wire multm_reduce_qs108;
  wire multm_reduce_qs109;
  wire multm_reduce_qs110;
  wire multm_reduce_qs111;
  wire multm_reduce_qs112;
  wire multm_reduce_qs113;
  wire multm_reduce_qs114;
  wire multm_reduce_qs115;
  wire multm_reduce_qs116;
  wire multm_reduce_qs117;
  wire multm_reduce_qs118;
  wire multm_reduce_qs119;
  wire multm_reduce_qs120;
  wire multm_reduce_qs121;
  wire multm_reduce_qs122;
  wire multm_reduce_qs123;
  wire multm_reduce_qs124;
  wire multm_reduce_qs125;
  wire multm_reduce_qs126;
  wire multm_reduce_qs127;
  wire multm_reduce_qs128;
  wire multm_reduce_qs129;
  wire multm_reduce_qs130;
  wire multm_reduce_qs131;
  wire multm_reduce_qs132;
  wire multm_reduce_qs133;
  wire multm_reduce_qs134;
  wire multm_reduce_qs135;
  wire multm_reduce_qs136;
  wire multm_reduce_qs137;
  wire multm_reduce_qs138;
  wire multm_reduce_qs139;
  wire multm_reduce_qs140;
  wire multm_reduce_qs141;
  wire multm_reduce_qs142;
  wire multm_reduce_qs143;
  wire multm_reduce_qs144;
  wire multm_reduce_qs145;
  wire multm_reduce_qs146;
  wire multm_reduce_qs147;
  wire multm_reduce_qs148;
  wire multm_reduce_qs149;
  wire multm_reduce_qs150;
  wire multm_reduce_qs151;
  wire multm_reduce_qs152;
  wire multm_reduce_qs153;
  wire multm_reduce_qs154;
  wire multm_reduce_qs155;
  wire multm_reduce_qs156;
  wire multm_reduce_qs157;
  wire multm_reduce_qs158;
  wire multm_reduce_qs159;
  wire multm_reduce_qs160;
  wire multm_reduce_qs161;
  wire multm_reduce_qs162;
  wire multm_reduce_qs163;
  wire multm_reduce_qs164;
  wire multm_reduce_qs165;
  wire multm_reduce_qs166;
  wire multm_reduce_qs167;
  wire multm_reduce_qs168;
  wire multm_reduce_qs169;
  wire multm_reduce_qs170;
  wire multm_reduce_qs171;
  wire multm_reduce_qs172;
  wire multm_reduce_qs173;
  wire multm_reduce_qs174;
  wire multm_reduce_qs175;
  wire multm_reduce_qs176;
  wire multm_reduce_qs177;
  wire multm_reduce_qs178;
  wire multm_reduce_qs179;
  wire multm_reduce_qs180;
  wire multm_reduce_qs181;
  wire multm_reduce_qs182;
  wire multm_reduce_qs183;
  wire multm_reduce_qs184;
  wire multm_reduce_sticky_q;
  wire multm_reduce_vb;
  wire multm_reduce_vc0;
  wire multm_reduce_vc1;
  wire multm_reduce_vc2;
  wire multm_reduce_vc3;
  wire multm_reduce_vc4;
  wire multm_reduce_vc5;
  wire multm_reduce_vc6;
  wire multm_reduce_vc7;
  wire multm_reduce_vc8;
  wire multm_reduce_vc9;
  wire multm_reduce_vc10;
  wire multm_reduce_vc11;
  wire multm_reduce_vc12;
  wire multm_reduce_vc13;
  wire multm_reduce_vc14;
  wire multm_reduce_vc15;
  wire multm_reduce_vc16;
  wire multm_reduce_vc17;
  wire multm_reduce_vc18;
  wire multm_reduce_vc19;
  wire multm_reduce_vc20;
  wire multm_reduce_vc21;
  wire multm_reduce_vc22;
  wire multm_reduce_vc23;
  wire multm_reduce_vc24;
  wire multm_reduce_vc25;
  wire multm_reduce_vc26;
  wire multm_reduce_vc27;
  wire multm_reduce_vc28;
  wire multm_reduce_vc29;
  wire multm_reduce_vc30;
  wire multm_reduce_vc31;
  wire multm_reduce_vc32;
  wire multm_reduce_vc33;
  wire multm_reduce_vc34;
  wire multm_reduce_vc35;
  wire multm_reduce_vc36;
  wire multm_reduce_vc37;
  wire multm_reduce_vc38;
  wire multm_reduce_vc39;
  wire multm_reduce_vc40;
  wire multm_reduce_vc41;
  wire multm_reduce_vc42;
  wire multm_reduce_vc43;
  wire multm_reduce_vc44;
  wire multm_reduce_vc45;
  wire multm_reduce_vc46;
  wire multm_reduce_vc47;
  wire multm_reduce_vc48;
  wire multm_reduce_vc49;
  wire multm_reduce_vc50;
  wire multm_reduce_vc51;
  wire multm_reduce_vc52;
  wire multm_reduce_vc53;
  wire multm_reduce_vc54;
  wire multm_reduce_vc55;
  wire multm_reduce_vc56;
  wire multm_reduce_vc57;
  wire multm_reduce_vc58;
  wire multm_reduce_vc59;
  wire multm_reduce_vc60;
  wire multm_reduce_vc61;
  wire multm_reduce_vc62;
  wire multm_reduce_vc63;
  wire multm_reduce_vc64;
  wire multm_reduce_vc65;
  wire multm_reduce_vc66;
  wire multm_reduce_vc67;
  wire multm_reduce_vc68;
  wire multm_reduce_vc69;
  wire multm_reduce_vc70;
  wire multm_reduce_vc71;
  wire multm_reduce_vc72;
  wire multm_reduce_vc73;
  wire multm_reduce_vc74;
  wire multm_reduce_vc75;
  wire multm_reduce_vc76;
  wire multm_reduce_vc77;
  wire multm_reduce_vc78;
  wire multm_reduce_vc79;
  wire multm_reduce_vc80;
  wire multm_reduce_vc81;
  wire multm_reduce_vc82;
  wire multm_reduce_vc83;
  wire multm_reduce_vc84;
  wire multm_reduce_vc85;
  wire multm_reduce_vc86;
  wire multm_reduce_vc87;
  wire multm_reduce_vc88;
  wire multm_reduce_vc89;
  wire multm_reduce_vc90;
  wire multm_reduce_vc91;
  wire multm_reduce_vc92;
  wire multm_reduce_vc93;
  wire multm_reduce_vc94;
  wire multm_reduce_vc95;
  wire multm_reduce_vc96;
  wire multm_reduce_vc97;
  wire multm_reduce_vc98;
  wire multm_reduce_vc99;
  wire multm_reduce_vc100;
  wire multm_reduce_vc101;
  wire multm_reduce_vc102;
  wire multm_reduce_vc103;
  wire multm_reduce_vc104;
  wire multm_reduce_vc105;
  wire multm_reduce_vc106;
  wire multm_reduce_vc107;
  wire multm_reduce_vc108;
  wire multm_reduce_vc109;
  wire multm_reduce_vc110;
  wire multm_reduce_vc111;
  wire multm_reduce_vc112;
  wire multm_reduce_vc113;
  wire multm_reduce_vc114;
  wire multm_reduce_vc115;
  wire multm_reduce_vc116;
  wire multm_reduce_vc117;
  wire multm_reduce_vc118;
  wire multm_reduce_vc119;
  wire multm_reduce_vc120;
  wire multm_reduce_vc121;
  wire multm_reduce_vc122;
  wire multm_reduce_vc123;
  wire multm_reduce_vc124;
  wire multm_reduce_vc125;
  wire multm_reduce_vc126;
  wire multm_reduce_vc127;
  wire multm_reduce_vc128;
  wire multm_reduce_vc129;
  wire multm_reduce_vc130;
  wire multm_reduce_vc131;
  wire multm_reduce_vc132;
  wire multm_reduce_vc133;
  wire multm_reduce_vc134;
  wire multm_reduce_vc135;
  wire multm_reduce_vc136;
  wire multm_reduce_vc137;
  wire multm_reduce_vc138;
  wire multm_reduce_vc139;
  wire multm_reduce_vc140;
  wire multm_reduce_vc141;
  wire multm_reduce_vc142;
  wire multm_reduce_vc143;
  wire multm_reduce_vc144;
  wire multm_reduce_vc145;
  wire multm_reduce_vc146;
  wire multm_reduce_vc147;
  wire multm_reduce_vc148;
  wire multm_reduce_vc149;
  wire multm_reduce_vc150;
  wire multm_reduce_vc151;
  wire multm_reduce_vc152;
  wire multm_reduce_vc153;
  wire multm_reduce_vc154;
  wire multm_reduce_vc155;
  wire multm_reduce_vc156;
  wire multm_reduce_vc157;
  wire multm_reduce_vc158;
  wire multm_reduce_vc159;
  wire multm_reduce_vc160;
  wire multm_reduce_vc161;
  wire multm_reduce_vc162;
  wire multm_reduce_vc163;
  wire multm_reduce_vc164;
  wire multm_reduce_vc165;
  wire multm_reduce_vc166;
  wire multm_reduce_vc167;
  wire multm_reduce_vc168;
  wire multm_reduce_vc169;
  wire multm_reduce_vc170;
  wire multm_reduce_vc171;
  wire multm_reduce_vc172;
  wire multm_reduce_vc173;
  wire multm_reduce_vc174;
  wire multm_reduce_vc175;
  wire multm_reduce_vc176;
  wire multm_reduce_vc177;
  wire multm_reduce_vc178;
  wire multm_reduce_vc179;
  wire multm_reduce_vc180;
  wire multm_reduce_vc181;
  wire multm_reduce_vc182;
  wire multm_reduce_vs0;
  wire multm_reduce_vs1;
  wire multm_reduce_vs2;
  wire multm_reduce_vs3;
  wire multm_reduce_vs4;
  wire multm_reduce_vs5;
  wire multm_reduce_vs6;
  wire multm_reduce_vs7;
  wire multm_reduce_vs8;
  wire multm_reduce_vs9;
  wire multm_reduce_vs10;
  wire multm_reduce_vs11;
  wire multm_reduce_vs12;
  wire multm_reduce_vs13;
  wire multm_reduce_vs14;
  wire multm_reduce_vs15;
  wire multm_reduce_vs16;
  wire multm_reduce_vs17;
  wire multm_reduce_vs18;
  wire multm_reduce_vs19;
  wire multm_reduce_vs20;
  wire multm_reduce_vs21;
  wire multm_reduce_vs22;
  wire multm_reduce_vs23;
  wire multm_reduce_vs24;
  wire multm_reduce_vs25;
  wire multm_reduce_vs26;
  wire multm_reduce_vs27;
  wire multm_reduce_vs28;
  wire multm_reduce_vs29;
  wire multm_reduce_vs30;
  wire multm_reduce_vs31;
  wire multm_reduce_vs32;
  wire multm_reduce_vs33;
  wire multm_reduce_vs34;
  wire multm_reduce_vs35;
  wire multm_reduce_vs36;
  wire multm_reduce_vs37;
  wire multm_reduce_vs38;
  wire multm_reduce_vs39;
  wire multm_reduce_vs40;
  wire multm_reduce_vs41;
  wire multm_reduce_vs42;
  wire multm_reduce_vs43;
  wire multm_reduce_vs44;
  wire multm_reduce_vs45;
  wire multm_reduce_vs46;
  wire multm_reduce_vs47;
  wire multm_reduce_vs48;
  wire multm_reduce_vs49;
  wire multm_reduce_vs50;
  wire multm_reduce_vs51;
  wire multm_reduce_vs52;
  wire multm_reduce_vs53;
  wire multm_reduce_vs54;
  wire multm_reduce_vs55;
  wire multm_reduce_vs56;
  wire multm_reduce_vs57;
  wire multm_reduce_vs58;
  wire multm_reduce_vs59;
  wire multm_reduce_vs60;
  wire multm_reduce_vs61;
  wire multm_reduce_vs62;
  wire multm_reduce_vs63;
  wire multm_reduce_vs64;
  wire multm_reduce_vs65;
  wire multm_reduce_vs66;
  wire multm_reduce_vs67;
  wire multm_reduce_vs68;
  wire multm_reduce_vs69;
  wire multm_reduce_vs70;
  wire multm_reduce_vs71;
  wire multm_reduce_vs72;
  wire multm_reduce_vs73;
  wire multm_reduce_vs74;
  wire multm_reduce_vs75;
  wire multm_reduce_vs76;
  wire multm_reduce_vs77;
  wire multm_reduce_vs78;
  wire multm_reduce_vs79;
  wire multm_reduce_vs80;
  wire multm_reduce_vs81;
  wire multm_reduce_vs82;
  wire multm_reduce_vs83;
  wire multm_reduce_vs84;
  wire multm_reduce_vs85;
  wire multm_reduce_vs86;
  wire multm_reduce_vs87;
  wire multm_reduce_vs88;
  wire multm_reduce_vs89;
  wire multm_reduce_vs90;
  wire multm_reduce_vs91;
  wire multm_reduce_vs92;
  wire multm_reduce_vs93;
  wire multm_reduce_vs94;
  wire multm_reduce_vs95;
  wire multm_reduce_vs96;
  wire multm_reduce_vs97;
  wire multm_reduce_vs98;
  wire multm_reduce_vs99;
  wire multm_reduce_vs100;
  wire multm_reduce_vs101;
  wire multm_reduce_vs102;
  wire multm_reduce_vs103;
  wire multm_reduce_vs104;
  wire multm_reduce_vs105;
  wire multm_reduce_vs106;
  wire multm_reduce_vs107;
  wire multm_reduce_vs108;
  wire multm_reduce_vs109;
  wire multm_reduce_vs110;
  wire multm_reduce_vs111;
  wire multm_reduce_vs112;
  wire multm_reduce_vs113;
  wire multm_reduce_vs114;
  wire multm_reduce_vs115;
  wire multm_reduce_vs116;
  wire multm_reduce_vs117;
  wire multm_reduce_vs118;
  wire multm_reduce_vs119;
  wire multm_reduce_vs120;
  wire multm_reduce_vs121;
  wire multm_reduce_vs122;
  wire multm_reduce_vs123;
  wire multm_reduce_vs124;
  wire multm_reduce_vs125;
  wire multm_reduce_vs126;
  wire multm_reduce_vs127;
  wire multm_reduce_vs128;
  wire multm_reduce_vs129;
  wire multm_reduce_vs130;
  wire multm_reduce_vs131;
  wire multm_reduce_vs132;
  wire multm_reduce_vs133;
  wire multm_reduce_vs134;
  wire multm_reduce_vs135;
  wire multm_reduce_vs136;
  wire multm_reduce_vs137;
  wire multm_reduce_vs138;
  wire multm_reduce_vs139;
  wire multm_reduce_vs140;
  wire multm_reduce_vs141;
  wire multm_reduce_vs142;
  wire multm_reduce_vs143;
  wire multm_reduce_vs144;
  wire multm_reduce_vs145;
  wire multm_reduce_vs146;
  wire multm_reduce_vs147;
  wire multm_reduce_vs148;
  wire multm_reduce_vs149;
  wire multm_reduce_vs150;
  wire multm_reduce_vs151;
  wire multm_reduce_vs152;
  wire multm_reduce_vs153;
  wire multm_reduce_vs154;
  wire multm_reduce_vs155;
  wire multm_reduce_vs156;
  wire multm_reduce_vs157;
  wire multm_reduce_vs158;
  wire multm_reduce_vs159;
  wire multm_reduce_vs160;
  wire multm_reduce_vs161;
  wire multm_reduce_vs162;
  wire multm_reduce_vs163;
  wire multm_reduce_vs164;
  wire multm_reduce_vs165;
  wire multm_reduce_vs166;
  wire multm_reduce_vs167;
  wire multm_reduce_vs168;
  wire multm_reduce_vs169;
  wire multm_reduce_vs170;
  wire multm_reduce_vs171;
  wire multm_reduce_vs172;
  wire multm_reduce_vs173;
  wire multm_reduce_vs174;
  wire multm_reduce_vs175;
  wire multm_reduce_vs176;
  wire multm_reduce_vs177;
  wire multm_reduce_vs178;
  wire multm_reduce_vs179;
  wire multm_reduce_vs180;
  wire multm_reduce_vs181;
  wire multm_reduce_vs182;
  wire multm_reduce_vt;
  wire nor2_zn;
  wire pcq0;
  wire pcq1;
  wire pcq2;
  wire pcq3;
  wire pcq4;
  wire pcq5;
  wire pcq6;
  wire pcq7;
  wire pcq8;
  wire pcq9;
  wire pcq10;
  wire pcq11;
  wire pcq12;
  wire pcq13;
  wire pcq14;
  wire pcq15;
  wire pcq16;
  wire pcq17;
  wire pcq18;
  wire pcq19;
  wire pcq20;
  wire pcq21;
  wire pcq22;
  wire pcq23;
  wire pcq24;
  wire pcq25;
  wire pcq26;
  wire pcq27;
  wire pcq28;
  wire pcq29;
  wire pcq30;
  wire pcq31;
  wire pcq32;
  wire pcq33;
  wire pcq34;
  wire pcq35;
  wire pcq36;
  wire pcq37;
  wire pcq38;
  wire pcq39;
  wire pcq40;
  wire pcq41;
  wire pcq42;
  wire pcq43;
  wire pcq44;
  wire pcq45;
  wire pcq46;
  wire pcq47;
  wire pcq48;
  wire pcq49;
  wire pcq50;
  wire pcq51;
  wire pcq52;
  wire pcq53;
  wire pcq54;
  wire pcq55;
  wire pcq56;
  wire pcq57;
  wire pcq58;
  wire pcq59;
  wire pcq60;
  wire pcq61;
  wire pcq62;
  wire pcq63;
  wire pcq64;
  wire pcq65;
  wire pcq66;
  wire pcq67;
  wire pcq68;
  wire pcq69;
  wire pcq70;
  wire pcq71;
  wire pcq72;
  wire pcq73;
  wire pcq74;
  wire pcq75;
  wire pcq76;
  wire pcq77;
  wire pcq78;
  wire pcq79;
  wire pcq80;
  wire pcq81;
  wire pcq82;
  wire pcq83;
  wire pcq84;
  wire pcq85;
  wire pcq86;
  wire pcq87;
  wire pcq88;
  wire pcq89;
  wire pcq90;
  wire pcq91;
  wire pcq92;
  wire pcq93;
  wire pcq94;
  wire pcq95;
  wire pcq96;
  wire pcq97;
  wire pcq98;
  wire pcq99;
  wire pcq100;
  wire pcq101;
  wire pcq102;
  wire pcq103;
  wire pcq104;
  wire pcq105;
  wire pcq106;
  wire pcq107;
  wire pcq108;
  wire pcq109;
  wire pcq110;
  wire pcq111;
  wire pcq112;
  wire pcq113;
  wire pcq114;
  wire pcq115;
  wire pcq116;
  wire pcq117;
  wire pcq118;
  wire pcq119;
  wire pcq120;
  wire pcq121;
  wire pcq122;
  wire pcq123;
  wire pcq124;
  wire pcq125;
  wire pcq126;
  wire pcq127;
  wire pcq128;
  wire pcq129;
  wire pcq130;
  wire pcq131;
  wire pcq132;
  wire pcq133;
  wire pcq134;
  wire pcq135;
  wire pcq136;
  wire pcq137;
  wire pcq138;
  wire pcq139;
  wire pcq140;
  wire pcq141;
  wire pcq142;
  wire pcq143;
  wire pcq144;
  wire pcq145;
  wire pcq146;
  wire pcq147;
  wire pcq148;
  wire pcq149;
  wire pcq150;
  wire pcq151;
  wire pcq152;
  wire pcq153;
  wire pcq154;
  wire pcq155;
  wire pcq156;
  wire pcq157;
  wire pcq158;
  wire pcq159;
  wire pcq160;
  wire pcq161;
  wire pcq162;
  wire pcq163;
  wire pcq164;
  wire pcq165;
  wire pcq166;
  wire pcq167;
  wire pcq168;
  wire pcq169;
  wire pcq170;
  wire pcq171;
  wire pcq172;
  wire pcq173;
  wire pcq174;
  wire pcq175;
  wire pcq176;
  wire pcq177;
  wire pcq178;
  wire pcq179;
  wire pcq180;
  wire pcq181;
  wire pcq182;
  wire pcq183;
  wire pcr0;
  wire pcr1;
  wire pcr2;
  wire pcr3;
  wire pcr4;
  wire pcr5;
  wire pcr6;
  wire pcr7;
  wire pcr8;
  wire pcr9;
  wire pcr10;
  wire pcr11;
  wire pcr12;
  wire pcr13;
  wire pcr14;
  wire pcr15;
  wire pcr16;
  wire pcr17;
  wire pcr18;
  wire pcr19;
  wire pcr20;
  wire pcr21;
  wire pcr22;
  wire pcr23;
  wire pcr24;
  wire pcr25;
  wire pcr26;
  wire pcr27;
  wire pcr28;
  wire pcr29;
  wire pcr30;
  wire pcr31;
  wire pcr32;
  wire pcr33;
  wire pcr34;
  wire pcr35;
  wire pcr36;
  wire pcr37;
  wire pcr38;
  wire pcr39;
  wire pcr40;
  wire pcr41;
  wire pcr42;
  wire pcr43;
  wire pcr44;
  wire pcr45;
  wire pcr46;
  wire pcr47;
  wire pcr48;
  wire pcr49;
  wire pcr50;
  wire pcr51;
  wire pcr52;
  wire pcr53;
  wire pcr54;
  wire pcr55;
  wire pcr56;
  wire pcr57;
  wire pcr58;
  wire pcr59;
  wire pcr60;
  wire pcr61;
  wire pcr62;
  wire pcr63;
  wire pcr64;
  wire pcr65;
  wire pcr66;
  wire pcr67;
  wire pcr68;
  wire pcr69;
  wire pcr70;
  wire pcr71;
  wire pcr72;
  wire pcr73;
  wire pcr74;
  wire pcr75;
  wire pcr76;
  wire pcr77;
  wire pcr78;
  wire pcr79;
  wire pcr80;
  wire pcr81;
  wire pcr82;
  wire pcr83;
  wire pcr84;
  wire pcr85;
  wire pcr86;
  wire pcr87;
  wire pcr88;
  wire pcr89;
  wire pcr90;
  wire pcr91;
  wire pcr92;
  wire pcr93;
  wire pcr94;
  wire pcr95;
  wire pcr96;
  wire pcr97;
  wire pcr98;
  wire pcr99;
  wire pcr100;
  wire pcr101;
  wire pcr102;
  wire pcr103;
  wire pcr104;
  wire pcr105;
  wire pcr106;
  wire pcr107;
  wire pcr108;
  wire pcr109;
  wire pcr110;
  wire pcr111;
  wire pcr112;
  wire pcr113;
  wire pcr114;
  wire pcr115;
  wire pcr116;
  wire pcr117;
  wire pcr118;
  wire pcr119;
  wire pcr120;
  wire pcr121;
  wire pcr122;
  wire pcr123;
  wire pcr124;
  wire pcr125;
  wire pcr126;
  wire pcr127;
  wire pcr128;
  wire pcr129;
  wire pcr130;
  wire pcr131;
  wire pcr132;
  wire pcr133;
  wire pcr134;
  wire pcr135;
  wire pcr136;
  wire pcr137;
  wire pcr138;
  wire pcr139;
  wire pcr140;
  wire pcr141;
  wire pcr142;
  wire pcr143;
  wire pcr144;
  wire pcr145;
  wire pcr146;
  wire pcr147;
  wire pcr148;
  wire pcr149;
  wire pcr150;
  wire pcr151;
  wire pcr152;
  wire pcr153;
  wire pcr154;
  wire pcr155;
  wire pcr156;
  wire pcr157;
  wire pcr158;
  wire pcr159;
  wire pcr160;
  wire pcr161;
  wire pcr162;
  wire pcr163;
  wire pcr164;
  wire pcr165;
  wire pcr166;
  wire pcr167;
  wire pcr168;
  wire pcr169;
  wire pcr170;
  wire pcr171;
  wire pcr172;
  wire pcr173;
  wire pcr174;
  wire pcr175;
  wire pcr176;
  wire pcr177;
  wire pcr178;
  wire pcr179;
  wire pcr180;
  wire pcr181;
  wire pcr182;
  wire pcr183;
  wire psq0;
  wire psq1;
  wire psq2;
  wire psq3;
  wire psq4;
  wire psq5;
  wire psq6;
  wire psq7;
  wire psq8;
  wire psq9;
  wire psq10;
  wire psq11;
  wire psq12;
  wire psq13;
  wire psq14;
  wire psq15;
  wire psq16;
  wire psq17;
  wire psq18;
  wire psq19;
  wire psq20;
  wire psq21;
  wire psq22;
  wire psq23;
  wire psq24;
  wire psq25;
  wire psq26;
  wire psq27;
  wire psq28;
  wire psq29;
  wire psq30;
  wire psq31;
  wire psq32;
  wire psq33;
  wire psq34;
  wire psq35;
  wire psq36;
  wire psq37;
  wire psq38;
  wire psq39;
  wire psq40;
  wire psq41;
  wire psq42;
  wire psq43;
  wire psq44;
  wire psq45;
  wire psq46;
  wire psq47;
  wire psq48;
  wire psq49;
  wire psq50;
  wire psq51;
  wire psq52;
  wire psq53;
  wire psq54;
  wire psq55;
  wire psq56;
  wire psq57;
  wire psq58;
  wire psq59;
  wire psq60;
  wire psq61;
  wire psq62;
  wire psq63;
  wire psq64;
  wire psq65;
  wire psq66;
  wire psq67;
  wire psq68;
  wire psq69;
  wire psq70;
  wire psq71;
  wire psq72;
  wire psq73;
  wire psq74;
  wire psq75;
  wire psq76;
  wire psq77;
  wire psq78;
  wire psq79;
  wire psq80;
  wire psq81;
  wire psq82;
  wire psq83;
  wire psq84;
  wire psq85;
  wire psq86;
  wire psq87;
  wire psq88;
  wire psq89;
  wire psq90;
  wire psq91;
  wire psq92;
  wire psq93;
  wire psq94;
  wire psq95;
  wire psq96;
  wire psq97;
  wire psq98;
  wire psq99;
  wire psq100;
  wire psq101;
  wire psq102;
  wire psq103;
  wire psq104;
  wire psq105;
  wire psq106;
  wire psq107;
  wire psq108;
  wire psq109;
  wire psq110;
  wire psq111;
  wire psq112;
  wire psq113;
  wire psq114;
  wire psq115;
  wire psq116;
  wire psq117;
  wire psq118;
  wire psq119;
  wire psq120;
  wire psq121;
  wire psq122;
  wire psq123;
  wire psq124;
  wire psq125;
  wire psq126;
  wire psq127;
  wire psq128;
  wire psq129;
  wire psq130;
  wire psq131;
  wire psq132;
  wire psq133;
  wire psq134;
  wire psq135;
  wire psq136;
  wire psq137;
  wire psq138;
  wire psq139;
  wire psq140;
  wire psq141;
  wire psq142;
  wire psq143;
  wire psq144;
  wire psq145;
  wire psq146;
  wire psq147;
  wire psq148;
  wire psq149;
  wire psq150;
  wire psq151;
  wire psq152;
  wire psq153;
  wire psq154;
  wire psq155;
  wire psq156;
  wire psq157;
  wire psq158;
  wire psq159;
  wire psq160;
  wire psq161;
  wire psq162;
  wire psq163;
  wire psq164;
  wire psq165;
  wire psq166;
  wire psq167;
  wire psq168;
  wire psq169;
  wire psq170;
  wire psq171;
  wire psq172;
  wire psq173;
  wire psq174;
  wire psq175;
  wire psq176;
  wire psq177;
  wire psq178;
  wire psq179;
  wire psq180;
  wire psq181;
  wire psq182;
  wire psq183;
  wire psr0;
  wire psr1;
  wire psr2;
  wire psr3;
  wire psr4;
  wire psr5;
  wire psr6;
  wire psr7;
  wire psr8;
  wire psr9;
  wire psr10;
  wire psr11;
  wire psr12;
  wire psr13;
  wire psr14;
  wire psr15;
  wire psr16;
  wire psr17;
  wire psr18;
  wire psr19;
  wire psr20;
  wire psr21;
  wire psr22;
  wire psr23;
  wire psr24;
  wire psr25;
  wire psr26;
  wire psr27;
  wire psr28;
  wire psr29;
  wire psr30;
  wire psr31;
  wire psr32;
  wire psr33;
  wire psr34;
  wire psr35;
  wire psr36;
  wire psr37;
  wire psr38;
  wire psr39;
  wire psr40;
  wire psr41;
  wire psr42;
  wire psr43;
  wire psr44;
  wire psr45;
  wire psr46;
  wire psr47;
  wire psr48;
  wire psr49;
  wire psr50;
  wire psr51;
  wire psr52;
  wire psr53;
  wire psr54;
  wire psr55;
  wire psr56;
  wire psr57;
  wire psr58;
  wire psr59;
  wire psr60;
  wire psr61;
  wire psr62;
  wire psr63;
  wire psr64;
  wire psr65;
  wire psr66;
  wire psr67;
  wire psr68;
  wire psr69;
  wire psr70;
  wire psr71;
  wire psr72;
  wire psr73;
  wire psr74;
  wire psr75;
  wire psr76;
  wire psr77;
  wire psr78;
  wire psr79;
  wire psr80;
  wire psr81;
  wire psr82;
  wire psr83;
  wire psr84;
  wire psr85;
  wire psr86;
  wire psr87;
  wire psr88;
  wire psr89;
  wire psr90;
  wire psr91;
  wire psr92;
  wire psr93;
  wire psr94;
  wire psr95;
  wire psr96;
  wire psr97;
  wire psr98;
  wire psr99;
  wire psr100;
  wire psr101;
  wire psr102;
  wire psr103;
  wire psr104;
  wire psr105;
  wire psr106;
  wire psr107;
  wire psr108;
  wire psr109;
  wire psr110;
  wire psr111;
  wire psr112;
  wire psr113;
  wire psr114;
  wire psr115;
  wire psr116;
  wire psr117;
  wire psr118;
  wire psr119;
  wire psr120;
  wire psr121;
  wire psr122;
  wire psr123;
  wire psr124;
  wire psr125;
  wire psr126;
  wire psr127;
  wire psr128;
  wire psr129;
  wire psr130;
  wire psr131;
  wire psr132;
  wire psr133;
  wire psr134;
  wire psr135;
  wire psr136;
  wire psr137;
  wire psr138;
  wire psr139;
  wire psr140;
  wire psr141;
  wire psr142;
  wire psr143;
  wire psr144;
  wire psr145;
  wire psr146;
  wire psr147;
  wire psr148;
  wire psr149;
  wire psr150;
  wire psr151;
  wire psr152;
  wire psr153;
  wire psr154;
  wire psr155;
  wire psr156;
  wire psr157;
  wire psr158;
  wire psr159;
  wire psr160;
  wire psr161;
  wire psr162;
  wire psr163;
  wire psr164;
  wire psr165;
  wire psr166;
  wire psr167;
  wire psr168;
  wire psr169;
  wire psr170;
  wire psr171;
  wire psr172;
  wire psr173;
  wire psr174;
  wire psr175;
  wire psr176;
  wire psr177;
  wire psr178;
  wire psr179;
  wire psr180;
  wire psr181;
  wire psr182;
  wire psr183;
  wire qc0;
  wire qc1;
  wire qc2;
  wire qc3;
  wire qc4;
  wire qc5;
  wire qc6;
  wire qc7;
  wire qc8;
  wire qc9;
  wire qc10;
  wire qc11;
  wire qc12;
  wire qc13;
  wire qc14;
  wire qc15;
  wire qc16;
  wire qc17;
  wire qc18;
  wire qc19;
  wire qc20;
  wire qc21;
  wire qc22;
  wire qc23;
  wire qc24;
  wire qc25;
  wire qc26;
  wire qc27;
  wire qc28;
  wire qc29;
  wire qc30;
  wire qc31;
  wire qc32;
  wire qc33;
  wire qc34;
  wire qc35;
  wire qc36;
  wire qc37;
  wire qc38;
  wire qc39;
  wire qc40;
  wire qc41;
  wire qc42;
  wire qc43;
  wire qc44;
  wire qc45;
  wire qc46;
  wire qc47;
  wire qc48;
  wire qc49;
  wire qc50;
  wire qc51;
  wire qc52;
  wire qc53;
  wire qc54;
  wire qc55;
  wire qc56;
  wire qc57;
  wire qc58;
  wire qc59;
  wire qc60;
  wire qc61;
  wire qc62;
  wire qc63;
  wire qc64;
  wire qc65;
  wire qc66;
  wire qc67;
  wire qc68;
  wire qc69;
  wire qc70;
  wire qc71;
  wire qc72;
  wire qc73;
  wire qc74;
  wire qc75;
  wire qc76;
  wire qc77;
  wire qc78;
  wire qc79;
  wire qc80;
  wire qc81;
  wire qc82;
  wire qc83;
  wire qc84;
  wire qc85;
  wire qc86;
  wire qc87;
  wire qc88;
  wire qc89;
  wire qc90;
  wire qc91;
  wire qc92;
  wire qc93;
  wire qc94;
  wire qc95;
  wire qc96;
  wire qc97;
  wire qc98;
  wire qc99;
  wire qc100;
  wire qc101;
  wire qc102;
  wire qc103;
  wire qc104;
  wire qc105;
  wire qc106;
  wire qc107;
  wire qc108;
  wire qc109;
  wire qc110;
  wire qc111;
  wire qc112;
  wire qc113;
  wire qc114;
  wire qc115;
  wire qc116;
  wire qc117;
  wire qc118;
  wire qc119;
  wire qc120;
  wire qc121;
  wire qc122;
  wire qc123;
  wire qc124;
  wire qc125;
  wire qc126;
  wire qc127;
  wire qc128;
  wire qc129;
  wire qc130;
  wire qc131;
  wire qc132;
  wire qc133;
  wire qc134;
  wire qc135;
  wire qc136;
  wire qc137;
  wire qc138;
  wire qc139;
  wire qc140;
  wire qc141;
  wire qc142;
  wire qc143;
  wire qc144;
  wire qc145;
  wire qc146;
  wire qc147;
  wire qc148;
  wire qc149;
  wire qc150;
  wire qc151;
  wire qc152;
  wire qc153;
  wire qc154;
  wire qc155;
  wire qc156;
  wire qc157;
  wire qc158;
  wire qc159;
  wire qc160;
  wire qc161;
  wire qc162;
  wire qc163;
  wire qc164;
  wire qc165;
  wire qc166;
  wire qc167;
  wire qc168;
  wire qc169;
  wire qc170;
  wire qc171;
  wire qc172;
  wire qc173;
  wire qc174;
  wire qc175;
  wire qc176;
  wire qc177;
  wire qc178;
  wire qc179;
  wire qc180;
  wire qc181;
  wire qc182;
  wire qc183;
  wire qs0;
  wire qs1;
  wire qs2;
  wire qs3;
  wire qs4;
  wire qs5;
  wire qs6;
  wire qs7;
  wire qs8;
  wire qs9;
  wire qs10;
  wire qs11;
  wire qs12;
  wire qs13;
  wire qs14;
  wire qs15;
  wire qs16;
  wire qs17;
  wire qs18;
  wire qs19;
  wire qs20;
  wire qs21;
  wire qs22;
  wire qs23;
  wire qs24;
  wire qs25;
  wire qs26;
  wire qs27;
  wire qs28;
  wire qs29;
  wire qs30;
  wire qs31;
  wire qs32;
  wire qs33;
  wire qs34;
  wire qs35;
  wire qs36;
  wire qs37;
  wire qs38;
  wire qs39;
  wire qs40;
  wire qs41;
  wire qs42;
  wire qs43;
  wire qs44;
  wire qs45;
  wire qs46;
  wire qs47;
  wire qs48;
  wire qs49;
  wire qs50;
  wire qs51;
  wire qs52;
  wire qs53;
  wire qs54;
  wire qs55;
  wire qs56;
  wire qs57;
  wire qs58;
  wire qs59;
  wire qs60;
  wire qs61;
  wire qs62;
  wire qs63;
  wire qs64;
  wire qs65;
  wire qs66;
  wire qs67;
  wire qs68;
  wire qs69;
  wire qs70;
  wire qs71;
  wire qs72;
  wire qs73;
  wire qs74;
  wire qs75;
  wire qs76;
  wire qs77;
  wire qs78;
  wire qs79;
  wire qs80;
  wire qs81;
  wire qs82;
  wire qs83;
  wire qs84;
  wire qs85;
  wire qs86;
  wire qs87;
  wire qs88;
  wire qs89;
  wire qs90;
  wire qs91;
  wire qs92;
  wire qs93;
  wire qs94;
  wire qs95;
  wire qs96;
  wire qs97;
  wire qs98;
  wire qs99;
  wire qs100;
  wire qs101;
  wire qs102;
  wire qs103;
  wire qs104;
  wire qs105;
  wire qs106;
  wire qs107;
  wire qs108;
  wire qs109;
  wire qs110;
  wire qs111;
  wire qs112;
  wire qs113;
  wire qs114;
  wire qs115;
  wire qs116;
  wire qs117;
  wire qs118;
  wire qs119;
  wire qs120;
  wire qs121;
  wire qs122;
  wire qs123;
  wire qs124;
  wire qs125;
  wire qs126;
  wire qs127;
  wire qs128;
  wire qs129;
  wire qs130;
  wire qs131;
  wire qs132;
  wire qs133;
  wire qs134;
  wire qs135;
  wire qs136;
  wire qs137;
  wire qs138;
  wire qs139;
  wire qs140;
  wire qs141;
  wire qs142;
  wire qs143;
  wire qs144;
  wire qs145;
  wire qs146;
  wire qs147;
  wire qs148;
  wire qs149;
  wire qs150;
  wire qs151;
  wire qs152;
  wire qs153;
  wire qs154;
  wire qs155;
  wire qs156;
  wire qs157;
  wire qs158;
  wire qs159;
  wire qs160;
  wire qs161;
  wire qs162;
  wire qs163;
  wire qs164;
  wire qs165;
  wire qs166;
  wire qs167;
  wire qs168;
  wire qs169;
  wire qs170;
  wire qs171;
  wire qs172;
  wire qs173;
  wire qs174;
  wire qs175;
  wire qs176;
  wire qs177;
  wire qs178;
  wire qs179;
  wire qs180;
  wire qs181;
  wire qs182;
  wire qs183;
  wire san;
  wire sap;
  wire saq;
  wire sar;
  wire sbp;
  wire sbq;
  wire sbr;
  wire srdd;
  wire xn0;
  wire xn1;
  wire xn2;
  wire xn3;
  wire xn4;
  wire xn5;
  wire xn6;

  assign ctre_cq0 = sadd & ctre_sp0;
  assign ctre_cq1 = ctre_sp1 & ctre_cp0;
  assign ctre_cq2 = ctre_sp2 & ctre_cp1;
  assign ctre_cq3 = ctre_sp3 & ctre_cp2;
  assign ctre_cq4 = ctre_sp4 & ctre_cp3;
  assign ctre_cq5 = ctre_sp5 & ctre_cp4;
  assign ctre_cq6 = ctre_sp6 & ctre_cp5;
  assign ctre_cq7 = ctre_sp7 & ctre_cp6;
  assign ctre_cq8 = ctre_sp8 & ctre_cp7;
  assign ctre_cq9 = ctre_sp9 & ctre_cp8;
  assign ctre_cr0 = xn5 & ctre_cq0;
  assign ctre_cr1 = xn5 & ctre_cq1;
  assign ctre_cr2 = xn5 & ctre_cq2;
  assign ctre_cr3 = xn5 & ctre_cq3;
  assign ctre_cr4 = xn5 & ctre_cq4;
  assign ctre_cr5 = xn5 & ctre_cq5;
  assign ctre_cr6 = xn5 & ctre_cq6;
  assign ctre_cr7 = xn5 & ctre_cq7;
  assign ctre_cr8 = xn5 & ctre_cq8;
  assign ctre_cr9 = xn5 & ctre_cq9;
  assign ctre_dq = ctre_dp | ctre_cp9;
  assign ctre_sq0 = sadd ^ ctre_sp0;
  assign ctre_sq1 = ctre_sp1 ^ ctre_cp0;
  assign ctre_sq2 = ctre_sp2 ^ ctre_cp1;
  assign ctre_sq3 = ctre_sp3 ^ ctre_cp2;
  assign ctre_sq4 = ctre_sp4 ^ ctre_cp3;
  assign ctre_sq5 = ctre_sp5 ^ ctre_cp4;
  assign ctre_sq6 = ctre_sp6 ^ ctre_cp5;
  assign ctre_sq7 = ctre_sp7 ^ ctre_cp6;
  assign ctre_sq8 = ctre_sp8 ^ ctre_cp7;
  assign ctre_sq9 = ctre_sp9 ^ ctre_cp8;
  assign ctre_sr0 = srdd | ctre_sq0;
  assign ctre_sr1 = xn5 & ctre_sq1;
  assign ctre_sr2 = xn5 & ctre_sq2;
  assign ctre_sr3 = srdd | ctre_sq3;
  assign ctre_sr4 = srdd | ctre_sq4;
  assign ctre_sr5 = xn5 & ctre_sq5;
  assign ctre_sr6 = xn5 & ctre_sq6;
  assign ctre_sr7 = xn5 & ctre_sq7;
  assign ctre_sr8 = xn5 & ctre_sq8;
  assign ctre_sr9 = xn5 & ctre_sq9;
  assign dn_o = ~nor2_zn;
  assign jp = multm_ctrp_ds & multm_ctrp_pulse_xn;
  assign jpn = ~jp;
  assign md = xn5 & ctre_dq;
  assign mdn = ~md;
  assign multm_compress_add3b_maj3b_or3b_wx0 = multm_compress_add3b_maj3b_wx0 | multm_compress_add3b_maj3b_wy0;
  assign multm_compress_add3b_maj3b_or3b_wx2 = multm_compress_add3b_maj3b_wx2 | multm_compress_add3b_maj3b_wy2;
  assign multm_compress_add3b_maj3b_or3b_wx3 = multm_compress_add3b_maj3b_wx3 | multm_compress_add3b_maj3b_wy3;
  assign multm_compress_add3b_maj3b_or3b_wx4 = multm_compress_add3b_maj3b_wx4 | multm_compress_add3b_maj3b_wy4;
  assign multm_compress_add3b_maj3b_or3b_wx5 = multm_compress_add3b_maj3b_wx5 | multm_compress_add3b_maj3b_wy5;
  assign multm_compress_add3b_maj3b_or3b_wx8 = multm_compress_add3b_maj3b_wx8 | multm_compress_add3b_maj3b_wy8;
  assign multm_compress_add3b_maj3b_or3b_wx9 = multm_compress_add3b_maj3b_wx9 | multm_compress_add3b_maj3b_wy9;
  assign multm_compress_add3b_maj3b_or3b_wx10 = multm_compress_add3b_maj3b_wx10 | multm_compress_add3b_maj3b_wy10;
  assign multm_compress_add3b_maj3b_or3b_wx11 = multm_compress_add3b_maj3b_wx11 | multm_compress_add3b_maj3b_wy11;
  assign multm_compress_add3b_maj3b_or3b_wx12 = multm_compress_add3b_maj3b_wx12 | multm_compress_add3b_maj3b_wy12;
  assign multm_compress_add3b_maj3b_or3b_wx13 = multm_compress_add3b_maj3b_wx13 | multm_compress_add3b_maj3b_wy13;
  assign multm_compress_add3b_maj3b_or3b_wx14 = multm_compress_add3b_maj3b_wx14 | multm_compress_add3b_maj3b_wy14;
  assign multm_compress_add3b_maj3b_or3b_wx15 = multm_compress_add3b_maj3b_wx15 | multm_compress_add3b_maj3b_wy15;
  assign multm_compress_add3b_maj3b_or3b_wx16 = multm_compress_add3b_maj3b_wx16 | multm_compress_add3b_maj3b_wy16;
  assign multm_compress_add3b_maj3b_or3b_wx17 = multm_compress_add3b_maj3b_wx17 | multm_compress_add3b_maj3b_wy17;
  assign multm_compress_add3b_maj3b_or3b_wx18 = multm_compress_add3b_maj3b_wx18 | multm_compress_add3b_maj3b_wy18;
  assign multm_compress_add3b_maj3b_or3b_wx19 = multm_compress_add3b_maj3b_wx19 | multm_compress_add3b_maj3b_wy19;
  assign multm_compress_add3b_maj3b_or3b_wx20 = multm_compress_add3b_maj3b_wx20 | multm_compress_add3b_maj3b_wy20;
  assign multm_compress_add3b_maj3b_or3b_wx21 = multm_compress_add3b_maj3b_wx21 | multm_compress_add3b_maj3b_wy21;
  assign multm_compress_add3b_maj3b_or3b_wx22 = multm_compress_add3b_maj3b_wx22 | multm_compress_add3b_maj3b_wy22;
  assign multm_compress_add3b_maj3b_or3b_wx23 = multm_compress_add3b_maj3b_wx23 | multm_compress_add3b_maj3b_wy23;
  assign multm_compress_add3b_maj3b_or3b_wx25 = multm_compress_add3b_maj3b_wx25 | multm_compress_add3b_maj3b_wy25;
  assign multm_compress_add3b_maj3b_or3b_wx26 = multm_compress_add3b_maj3b_wx26 | multm_compress_add3b_maj3b_wy26;
  assign multm_compress_add3b_maj3b_or3b_wx27 = multm_compress_add3b_maj3b_wx27 | multm_compress_add3b_maj3b_wy27;
  assign multm_compress_add3b_maj3b_or3b_wx28 = multm_compress_add3b_maj3b_wx28 | multm_compress_add3b_maj3b_wy28;
  assign multm_compress_add3b_maj3b_or3b_wx29 = multm_compress_add3b_maj3b_wx29 | multm_compress_add3b_maj3b_wy29;
  assign multm_compress_add3b_maj3b_or3b_wx30 = multm_compress_add3b_maj3b_wx30 | multm_compress_add3b_maj3b_wy30;
  assign multm_compress_add3b_maj3b_or3b_wx31 = multm_compress_add3b_maj3b_wx31 | multm_compress_add3b_maj3b_wy31;
  assign multm_compress_add3b_maj3b_or3b_wx32 = multm_compress_add3b_maj3b_wx32 | multm_compress_add3b_maj3b_wy32;
  assign multm_compress_add3b_maj3b_or3b_wx33 = multm_compress_add3b_maj3b_wx33 | multm_compress_add3b_maj3b_wy33;
  assign multm_compress_add3b_maj3b_or3b_wx34 = multm_compress_add3b_maj3b_wx34 | multm_compress_add3b_maj3b_wy34;
  assign multm_compress_add3b_maj3b_or3b_wx35 = multm_compress_add3b_maj3b_wx35 | multm_compress_add3b_maj3b_wy35;
  assign multm_compress_add3b_maj3b_or3b_wx36 = multm_compress_add3b_maj3b_wx36 | multm_compress_add3b_maj3b_wy36;
  assign multm_compress_add3b_maj3b_or3b_wx37 = multm_compress_add3b_maj3b_wx37 | multm_compress_add3b_maj3b_wy37;
  assign multm_compress_add3b_maj3b_or3b_wx38 = multm_compress_add3b_maj3b_wx38 | multm_compress_add3b_maj3b_wy38;
  assign multm_compress_add3b_maj3b_or3b_wx39 = multm_compress_add3b_maj3b_wx39 | multm_compress_add3b_maj3b_wy39;
  assign multm_compress_add3b_maj3b_or3b_wx40 = multm_compress_add3b_maj3b_wx40 | multm_compress_add3b_maj3b_wy40;
  assign multm_compress_add3b_maj3b_or3b_wx41 = multm_compress_add3b_maj3b_wx41 | multm_compress_add3b_maj3b_wy41;
  assign multm_compress_add3b_maj3b_or3b_wx44 = multm_compress_add3b_maj3b_wx44 | multm_compress_add3b_maj3b_wy44;
  assign multm_compress_add3b_maj3b_or3b_wx45 = multm_compress_add3b_maj3b_wx45 | multm_compress_add3b_maj3b_wy45;
  assign multm_compress_add3b_maj3b_or3b_wx46 = multm_compress_add3b_maj3b_wx46 | multm_compress_add3b_maj3b_wy46;
  assign multm_compress_add3b_maj3b_or3b_wx47 = multm_compress_add3b_maj3b_wx47 | multm_compress_add3b_maj3b_wy47;
  assign multm_compress_add3b_maj3b_or3b_wx48 = multm_compress_add3b_maj3b_wx48 | multm_compress_add3b_maj3b_wy48;
  assign multm_compress_add3b_maj3b_or3b_wx49 = multm_compress_add3b_maj3b_wx49 | multm_compress_add3b_maj3b_wy49;
  assign multm_compress_add3b_maj3b_or3b_wx50 = multm_compress_add3b_maj3b_wx50 | multm_compress_add3b_maj3b_wy50;
  assign multm_compress_add3b_maj3b_or3b_wx51 = multm_compress_add3b_maj3b_wx51 | multm_compress_add3b_maj3b_wy51;
  assign multm_compress_add3b_maj3b_or3b_wx52 = multm_compress_add3b_maj3b_wx52 | multm_compress_add3b_maj3b_wy52;
  assign multm_compress_add3b_maj3b_or3b_wx56 = multm_compress_add3b_maj3b_wx56 | multm_compress_add3b_maj3b_wy56;
  assign multm_compress_add3b_maj3b_or3b_wx57 = multm_compress_add3b_maj3b_wx57 | multm_compress_add3b_maj3b_wy57;
  assign multm_compress_add3b_maj3b_or3b_wx58 = multm_compress_add3b_maj3b_wx58 | multm_compress_add3b_maj3b_wy58;
  assign multm_compress_add3b_maj3b_or3b_wx59 = multm_compress_add3b_maj3b_wx59 | multm_compress_add3b_maj3b_wy59;
  assign multm_compress_add3b_maj3b_or3b_wx60 = multm_compress_add3b_maj3b_wx60 | multm_compress_add3b_maj3b_wy60;
  assign multm_compress_add3b_maj3b_or3b_wx61 = multm_compress_add3b_maj3b_wx61 | multm_compress_add3b_maj3b_wy61;
  assign multm_compress_add3b_maj3b_or3b_wx62 = multm_compress_add3b_maj3b_wx62 | multm_compress_add3b_maj3b_wy62;
  assign multm_compress_add3b_maj3b_or3b_wx63 = multm_compress_add3b_maj3b_wx63 | multm_compress_add3b_maj3b_wy63;
  assign multm_compress_add3b_maj3b_or3b_wx64 = multm_compress_add3b_maj3b_wx64 | multm_compress_add3b_maj3b_wy64;
  assign multm_compress_add3b_maj3b_or3b_wx65 = multm_compress_add3b_maj3b_wx65 | multm_compress_add3b_maj3b_wy65;
  assign multm_compress_add3b_maj3b_or3b_wx66 = multm_compress_add3b_maj3b_wx66 | multm_compress_add3b_maj3b_wy66;
  assign multm_compress_add3b_maj3b_or3b_wx67 = multm_compress_add3b_maj3b_wx67 | multm_compress_add3b_maj3b_wy67;
  assign multm_compress_add3b_maj3b_or3b_wx68 = multm_compress_add3b_maj3b_wx68 | multm_compress_add3b_maj3b_wy68;
  assign multm_compress_add3b_maj3b_or3b_wx69 = multm_compress_add3b_maj3b_wx69 | multm_compress_add3b_maj3b_wy69;
  assign multm_compress_add3b_maj3b_or3b_wx70 = multm_compress_add3b_maj3b_wx70 | multm_compress_add3b_maj3b_wy70;
  assign multm_compress_add3b_maj3b_or3b_wx71 = multm_compress_add3b_maj3b_wx71 | multm_compress_add3b_maj3b_wy71;
  assign multm_compress_add3b_maj3b_or3b_wx72 = multm_compress_add3b_maj3b_wx72 | multm_compress_add3b_maj3b_wy72;
  assign multm_compress_add3b_maj3b_or3b_wx73 = multm_compress_add3b_maj3b_wx73 | multm_compress_add3b_maj3b_wy73;
  assign multm_compress_add3b_maj3b_or3b_wx75 = multm_compress_add3b_maj3b_wx75 | multm_compress_add3b_maj3b_wy75;
  assign multm_compress_add3b_maj3b_or3b_wx76 = multm_compress_add3b_maj3b_wx76 | multm_compress_add3b_maj3b_wy76;
  assign multm_compress_add3b_maj3b_or3b_wx77 = multm_compress_add3b_maj3b_wx77 | multm_compress_add3b_maj3b_wy77;
  assign multm_compress_add3b_maj3b_or3b_wx78 = multm_compress_add3b_maj3b_wx78 | multm_compress_add3b_maj3b_wy78;
  assign multm_compress_add3b_maj3b_or3b_wx79 = multm_compress_add3b_maj3b_wx79 | multm_compress_add3b_maj3b_wy79;
  assign multm_compress_add3b_maj3b_or3b_wx80 = multm_compress_add3b_maj3b_wx80 | multm_compress_add3b_maj3b_wy80;
  assign multm_compress_add3b_maj3b_or3b_wx81 = multm_compress_add3b_maj3b_wx81 | multm_compress_add3b_maj3b_wy81;
  assign multm_compress_add3b_maj3b_or3b_wx82 = multm_compress_add3b_maj3b_wx82 | multm_compress_add3b_maj3b_wy82;
  assign multm_compress_add3b_maj3b_or3b_wx83 = multm_compress_add3b_maj3b_wx83 | multm_compress_add3b_maj3b_wy83;
  assign multm_compress_add3b_maj3b_or3b_wx84 = multm_compress_add3b_maj3b_wx84 | multm_compress_add3b_maj3b_wy84;
  assign multm_compress_add3b_maj3b_or3b_wx85 = multm_compress_add3b_maj3b_wx85 | multm_compress_add3b_maj3b_wy85;
  assign multm_compress_add3b_maj3b_or3b_wx86 = multm_compress_add3b_maj3b_wx86 | multm_compress_add3b_maj3b_wy86;
  assign multm_compress_add3b_maj3b_or3b_wx87 = multm_compress_add3b_maj3b_wx87 | multm_compress_add3b_maj3b_wy87;
  assign multm_compress_add3b_maj3b_or3b_wx88 = multm_compress_add3b_maj3b_wx88 | multm_compress_add3b_maj3b_wy88;
  assign multm_compress_add3b_maj3b_or3b_wx89 = multm_compress_add3b_maj3b_wx89 | multm_compress_add3b_maj3b_wy89;
  assign multm_compress_add3b_maj3b_or3b_wx90 = multm_compress_add3b_maj3b_wx90 | multm_compress_add3b_maj3b_wy90;
  assign multm_compress_add3b_maj3b_or3b_wx91 = multm_compress_add3b_maj3b_wx91 | multm_compress_add3b_maj3b_wy91;
  assign multm_compress_add3b_maj3b_or3b_wx92 = multm_compress_add3b_maj3b_wx92 | multm_compress_add3b_maj3b_wy92;
  assign multm_compress_add3b_maj3b_or3b_wx93 = multm_compress_add3b_maj3b_wx93 | multm_compress_add3b_maj3b_wy93;
  assign multm_compress_add3b_maj3b_or3b_wx94 = multm_compress_add3b_maj3b_wx94 | multm_compress_add3b_maj3b_wy94;
  assign multm_compress_add3b_maj3b_or3b_wx95 = multm_compress_add3b_maj3b_wx95 | multm_compress_add3b_maj3b_wy95;
  assign multm_compress_add3b_maj3b_or3b_wx96 = multm_compress_add3b_maj3b_wx96 | multm_compress_add3b_maj3b_wy96;
  assign multm_compress_add3b_maj3b_or3b_wx97 = multm_compress_add3b_maj3b_wx97 | multm_compress_add3b_maj3b_wy97;
  assign multm_compress_add3b_maj3b_or3b_wx98 = multm_compress_add3b_maj3b_wx98 | multm_compress_add3b_maj3b_wy98;
  assign multm_compress_add3b_maj3b_or3b_wx99 = multm_compress_add3b_maj3b_wx99 | multm_compress_add3b_maj3b_wy99;
  assign multm_compress_add3b_maj3b_or3b_wx100 = multm_compress_add3b_maj3b_wx100 | multm_compress_add3b_maj3b_wy100;
  assign multm_compress_add3b_maj3b_or3b_wx103 = multm_compress_add3b_maj3b_wx103 | multm_compress_add3b_maj3b_wy103;
  assign multm_compress_add3b_maj3b_or3b_wx104 = multm_compress_add3b_maj3b_wx104 | multm_compress_add3b_maj3b_wy104;
  assign multm_compress_add3b_maj3b_or3b_wx106 = multm_compress_add3b_maj3b_wx106 | multm_compress_add3b_maj3b_wy106;
  assign multm_compress_add3b_maj3b_or3b_wx107 = multm_compress_add3b_maj3b_wx107 | multm_compress_add3b_maj3b_wy107;
  assign multm_compress_add3b_maj3b_or3b_wx111 = multm_compress_add3b_maj3b_wx111 | multm_compress_add3b_maj3b_wy111;
  assign multm_compress_add3b_maj3b_or3b_wx112 = multm_compress_add3b_maj3b_wx112 | multm_compress_add3b_maj3b_wy112;
  assign multm_compress_add3b_maj3b_or3b_wx113 = multm_compress_add3b_maj3b_wx113 | multm_compress_add3b_maj3b_wy113;
  assign multm_compress_add3b_maj3b_or3b_wx114 = multm_compress_add3b_maj3b_wx114 | multm_compress_add3b_maj3b_wy114;
  assign multm_compress_add3b_maj3b_or3b_wx115 = multm_compress_add3b_maj3b_wx115 | multm_compress_add3b_maj3b_wy115;
  assign multm_compress_add3b_maj3b_or3b_wx116 = multm_compress_add3b_maj3b_wx116 | multm_compress_add3b_maj3b_wy116;
  assign multm_compress_add3b_maj3b_or3b_wx117 = multm_compress_add3b_maj3b_wx117 | multm_compress_add3b_maj3b_wy117;
  assign multm_compress_add3b_maj3b_or3b_wx118 = multm_compress_add3b_maj3b_wx118 | multm_compress_add3b_maj3b_wy118;
  assign multm_compress_add3b_maj3b_or3b_wx124 = multm_compress_add3b_maj3b_wx124 | multm_compress_add3b_maj3b_wy124;
  assign multm_compress_add3b_maj3b_or3b_wx125 = multm_compress_add3b_maj3b_wx125 | multm_compress_add3b_maj3b_wy125;
  assign multm_compress_add3b_maj3b_or3b_wx126 = multm_compress_add3b_maj3b_wx126 | multm_compress_add3b_maj3b_wy126;
  assign multm_compress_add3b_maj3b_or3b_wx127 = multm_compress_add3b_maj3b_wx127 | multm_compress_add3b_maj3b_wy127;
  assign multm_compress_add3b_maj3b_or3b_wx128 = multm_compress_add3b_maj3b_wx128 | multm_compress_add3b_maj3b_wy128;
  assign multm_compress_add3b_maj3b_or3b_wx129 = multm_compress_add3b_maj3b_wx129 | multm_compress_add3b_maj3b_wy129;
  assign multm_compress_add3b_maj3b_or3b_wx130 = multm_compress_add3b_maj3b_wx130 | multm_compress_add3b_maj3b_wy130;
  assign multm_compress_add3b_maj3b_or3b_wx131 = multm_compress_add3b_maj3b_wx131 | multm_compress_add3b_maj3b_wy131;
  assign multm_compress_add3b_maj3b_or3b_wx132 = multm_compress_add3b_maj3b_wx132 | multm_compress_add3b_maj3b_wy132;
  assign multm_compress_add3b_maj3b_or3b_wx133 = multm_compress_add3b_maj3b_wx133 | multm_compress_add3b_maj3b_wy133;
  assign multm_compress_add3b_maj3b_or3b_wx134 = multm_compress_add3b_maj3b_wx134 | multm_compress_add3b_maj3b_wy134;
  assign multm_compress_add3b_maj3b_or3b_wx135 = multm_compress_add3b_maj3b_wx135 | multm_compress_add3b_maj3b_wy135;
  assign multm_compress_add3b_maj3b_or3b_wx136 = multm_compress_add3b_maj3b_wx136 | multm_compress_add3b_maj3b_wy136;
  assign multm_compress_add3b_maj3b_or3b_wx137 = multm_compress_add3b_maj3b_wx137 | multm_compress_add3b_maj3b_wy137;
  assign multm_compress_add3b_maj3b_or3b_wx138 = multm_compress_add3b_maj3b_wx138 | multm_compress_add3b_maj3b_wy138;
  assign multm_compress_add3b_maj3b_or3b_wx139 = multm_compress_add3b_maj3b_wx139 | multm_compress_add3b_maj3b_wy139;
  assign multm_compress_add3b_maj3b_or3b_wx140 = multm_compress_add3b_maj3b_wx140 | multm_compress_add3b_maj3b_wy140;
  assign multm_compress_add3b_maj3b_or3b_wx141 = multm_compress_add3b_maj3b_wx141 | multm_compress_add3b_maj3b_wy141;
  assign multm_compress_add3b_maj3b_or3b_wx145 = multm_compress_add3b_maj3b_wx145 | multm_compress_add3b_maj3b_wy145;
  assign multm_compress_add3b_maj3b_or3b_wx146 = multm_compress_add3b_maj3b_wx146 | multm_compress_add3b_maj3b_wy146;
  assign multm_compress_add3b_maj3b_or3b_wx147 = multm_compress_add3b_maj3b_wx147 | multm_compress_add3b_maj3b_wy147;
  assign multm_compress_add3b_maj3b_or3b_wx148 = multm_compress_add3b_maj3b_wx148 | multm_compress_add3b_maj3b_wy148;
  assign multm_compress_add3b_maj3b_or3b_wx149 = multm_compress_add3b_maj3b_wx149 | multm_compress_add3b_maj3b_wy149;
  assign multm_compress_add3b_maj3b_or3b_wx150 = multm_compress_add3b_maj3b_wx150 | multm_compress_add3b_maj3b_wy150;
  assign multm_compress_add3b_maj3b_or3b_wx151 = multm_compress_add3b_maj3b_wx151 | multm_compress_add3b_maj3b_wy151;
  assign multm_compress_add3b_maj3b_or3b_wx154 = multm_compress_add3b_maj3b_wx154 | multm_compress_add3b_maj3b_wy154;
  assign multm_compress_add3b_maj3b_or3b_wx155 = multm_compress_add3b_maj3b_wx155 | multm_compress_add3b_maj3b_wy155;
  assign multm_compress_add3b_maj3b_or3b_wx161 = multm_compress_add3b_maj3b_wx161 | multm_compress_add3b_maj3b_wy161;
  assign multm_compress_add3b_maj3b_or3b_wx162 = multm_compress_add3b_maj3b_wx162 | multm_compress_add3b_maj3b_wy162;
  assign multm_compress_add3b_maj3b_or3b_wx163 = multm_compress_add3b_maj3b_wx163 | multm_compress_add3b_maj3b_wy163;
  assign multm_compress_add3b_maj3b_or3b_wx164 = multm_compress_add3b_maj3b_wx164 | multm_compress_add3b_maj3b_wy164;
  assign multm_compress_add3b_maj3b_or3b_wx165 = multm_compress_add3b_maj3b_wx165 | multm_compress_add3b_maj3b_wy165;
  assign multm_compress_add3b_maj3b_or3b_wx166 = multm_compress_add3b_maj3b_wx166 | multm_compress_add3b_maj3b_wy166;
  assign multm_compress_add3b_maj3b_or3b_wx167 = multm_compress_add3b_maj3b_wx167 | multm_compress_add3b_maj3b_wy167;
  assign multm_compress_add3b_maj3b_or3b_wx168 = multm_compress_add3b_maj3b_wx168 | multm_compress_add3b_maj3b_wy168;
  assign multm_compress_add3b_maj3b_or3b_wx169 = multm_compress_add3b_maj3b_wx169 | multm_compress_add3b_maj3b_wy169;
  assign multm_compress_add3b_maj3b_or3b_wx170 = multm_compress_add3b_maj3b_wx170 | multm_compress_add3b_maj3b_wy170;
  assign multm_compress_add3b_maj3b_or3b_wx171 = multm_compress_add3b_maj3b_wx171 | multm_compress_add3b_maj3b_wy171;
  assign multm_compress_add3b_maj3b_or3b_wx172 = multm_compress_add3b_maj3b_wx172 | multm_compress_add3b_maj3b_wy172;
  assign multm_compress_add3b_maj3b_or3b_wx176 = multm_compress_add3b_maj3b_wx176 | multm_compress_add3b_maj3b_wy176;
  assign multm_compress_add3b_maj3b_or3b_wx177 = multm_compress_add3b_maj3b_wx177 | multm_compress_add3b_maj3b_wy177;
  assign multm_compress_add3b_maj3b_or3b_wx178 = multm_compress_add3b_maj3b_wx178 | multm_compress_add3b_maj3b_wy178;
  assign multm_compress_add3b_maj3b_or3b_wx179 = multm_compress_add3b_maj3b_wx179 | multm_compress_add3b_maj3b_wy179;
  assign multm_compress_add3b_maj3b_or3b_wx180 = multm_compress_add3b_maj3b_wx180 | multm_compress_add3b_maj3b_wy180;
  assign multm_compress_add3b_maj3b_or3b_wx181 = multm_compress_add3b_maj3b_wx181 | multm_compress_add3b_maj3b_wy181;
  assign multm_compress_add3b_maj3b_or3b_wx182 = multm_compress_add3b_maj3b_wx182 | multm_compress_add3b_maj3b_wy182;
  assign multm_compress_add3b_maj3b_wx0 = multm_qsp1 & multm_qcp0;
  assign multm_compress_add3b_maj3b_wx2 = multm_qsp3 & multm_qcp2;
  assign multm_compress_add3b_maj3b_wx3 = multm_qsp4 & multm_qcp3;
  assign multm_compress_add3b_maj3b_wx4 = multm_qsp5 & multm_qcp4;
  assign multm_compress_add3b_maj3b_wx5 = multm_qsp6 & multm_qcp5;
  assign multm_compress_add3b_maj3b_wx8 = multm_qsp9 & multm_qcp8;
  assign multm_compress_add3b_maj3b_wx9 = multm_qsp10 & multm_qcp9;
  assign multm_compress_add3b_maj3b_wx10 = multm_qsp11 & multm_qcp10;
  assign multm_compress_add3b_maj3b_wx11 = multm_qsp12 & multm_qcp11;
  assign multm_compress_add3b_maj3b_wx12 = multm_qsp13 & multm_qcp12;
  assign multm_compress_add3b_maj3b_wx13 = multm_qsp14 & multm_qcp13;
  assign multm_compress_add3b_maj3b_wx14 = multm_qsp15 & multm_qcp14;
  assign multm_compress_add3b_maj3b_wx15 = multm_qsp16 & multm_qcp15;
  assign multm_compress_add3b_maj3b_wx16 = multm_qsp17 & multm_qcp16;
  assign multm_compress_add3b_maj3b_wx17 = multm_qsp18 & multm_qcp17;
  assign multm_compress_add3b_maj3b_wx18 = multm_qsp19 & multm_qcp18;
  assign multm_compress_add3b_maj3b_wx19 = multm_qsp20 & multm_qcp19;
  assign multm_compress_add3b_maj3b_wx20 = multm_qsp21 & multm_qcp20;
  assign multm_compress_add3b_maj3b_wx21 = multm_qsp22 & multm_qcp21;
  assign multm_compress_add3b_maj3b_wx22 = multm_qsp23 & multm_qcp22;
  assign multm_compress_add3b_maj3b_wx23 = multm_qsp24 & multm_qcp23;
  assign multm_compress_add3b_maj3b_wx25 = multm_qsp26 & multm_qcp25;
  assign multm_compress_add3b_maj3b_wx26 = multm_qsp27 & multm_qcp26;
  assign multm_compress_add3b_maj3b_wx27 = multm_qsp28 & multm_qcp27;
  assign multm_compress_add3b_maj3b_wx28 = multm_qsp29 & multm_qcp28;
  assign multm_compress_add3b_maj3b_wx29 = multm_qsp30 & multm_qcp29;
  assign multm_compress_add3b_maj3b_wx30 = multm_qsp31 & multm_qcp30;
  assign multm_compress_add3b_maj3b_wx31 = multm_qsp32 & multm_qcp31;
  assign multm_compress_add3b_maj3b_wx32 = multm_qsp33 & multm_qcp32;
  assign multm_compress_add3b_maj3b_wx33 = multm_qsp34 & multm_qcp33;
  assign multm_compress_add3b_maj3b_wx34 = multm_qsp35 & multm_qcp34;
  assign multm_compress_add3b_maj3b_wx35 = multm_qsp36 & multm_qcp35;
  assign multm_compress_add3b_maj3b_wx36 = multm_qsp37 & multm_qcp36;
  assign multm_compress_add3b_maj3b_wx37 = multm_qsp38 & multm_qcp37;
  assign multm_compress_add3b_maj3b_wx38 = multm_qsp39 & multm_qcp38;
  assign multm_compress_add3b_maj3b_wx39 = multm_qsp40 & multm_qcp39;
  assign multm_compress_add3b_maj3b_wx40 = multm_qsp41 & multm_qcp40;
  assign multm_compress_add3b_maj3b_wx41 = multm_qsp42 & multm_qcp41;
  assign multm_compress_add3b_maj3b_wx44 = multm_qsp45 & multm_qcp44;
  assign multm_compress_add3b_maj3b_wx45 = multm_qsp46 & multm_qcp45;
  assign multm_compress_add3b_maj3b_wx46 = multm_qsp47 & multm_qcp46;
  assign multm_compress_add3b_maj3b_wx47 = multm_qsp48 & multm_qcp47;
  assign multm_compress_add3b_maj3b_wx48 = multm_qsp49 & multm_qcp48;
  assign multm_compress_add3b_maj3b_wx49 = multm_qsp50 & multm_qcp49;
  assign multm_compress_add3b_maj3b_wx50 = multm_qsp51 & multm_qcp50;
  assign multm_compress_add3b_maj3b_wx51 = multm_qsp52 & multm_qcp51;
  assign multm_compress_add3b_maj3b_wx52 = multm_qsp53 & multm_qcp52;
  assign multm_compress_add3b_maj3b_wx56 = multm_qsp57 & multm_qcp56;
  assign multm_compress_add3b_maj3b_wx57 = multm_qsp58 & multm_qcp57;
  assign multm_compress_add3b_maj3b_wx58 = multm_qsp59 & multm_qcp58;
  assign multm_compress_add3b_maj3b_wx59 = multm_qsp60 & multm_qcp59;
  assign multm_compress_add3b_maj3b_wx60 = multm_qsp61 & multm_qcp60;
  assign multm_compress_add3b_maj3b_wx61 = multm_qsp62 & multm_qcp61;
  assign multm_compress_add3b_maj3b_wx62 = multm_qsp63 & multm_qcp62;
  assign multm_compress_add3b_maj3b_wx63 = multm_qsp64 & multm_qcp63;
  assign multm_compress_add3b_maj3b_wx64 = multm_qsp65 & multm_qcp64;
  assign multm_compress_add3b_maj3b_wx65 = multm_qsp66 & multm_qcp65;
  assign multm_compress_add3b_maj3b_wx66 = multm_qsp67 & multm_qcp66;
  assign multm_compress_add3b_maj3b_wx67 = multm_qsp68 & multm_qcp67;
  assign multm_compress_add3b_maj3b_wx68 = multm_qsp69 & multm_qcp68;
  assign multm_compress_add3b_maj3b_wx69 = multm_qsp70 & multm_qcp69;
  assign multm_compress_add3b_maj3b_wx70 = multm_qsp71 & multm_qcp70;
  assign multm_compress_add3b_maj3b_wx71 = multm_qsp72 & multm_qcp71;
  assign multm_compress_add3b_maj3b_wx72 = multm_qsp73 & multm_qcp72;
  assign multm_compress_add3b_maj3b_wx73 = multm_qsp74 & multm_qcp73;
  assign multm_compress_add3b_maj3b_wx75 = multm_qsp76 & multm_qcp75;
  assign multm_compress_add3b_maj3b_wx76 = multm_qsp77 & multm_qcp76;
  assign multm_compress_add3b_maj3b_wx77 = multm_qsp78 & multm_qcp77;
  assign multm_compress_add3b_maj3b_wx78 = multm_qsp79 & multm_qcp78;
  assign multm_compress_add3b_maj3b_wx79 = multm_qsp80 & multm_qcp79;
  assign multm_compress_add3b_maj3b_wx80 = multm_qsp81 & multm_qcp80;
  assign multm_compress_add3b_maj3b_wx81 = multm_qsp82 & multm_qcp81;
  assign multm_compress_add3b_maj3b_wx82 = multm_qsp83 & multm_qcp82;
  assign multm_compress_add3b_maj3b_wx83 = multm_qsp84 & multm_qcp83;
  assign multm_compress_add3b_maj3b_wx84 = multm_qsp85 & multm_qcp84;
  assign multm_compress_add3b_maj3b_wx85 = multm_qsp86 & multm_qcp85;
  assign multm_compress_add3b_maj3b_wx86 = multm_qsp87 & multm_qcp86;
  assign multm_compress_add3b_maj3b_wx87 = multm_qsp88 & multm_qcp87;
  assign multm_compress_add3b_maj3b_wx88 = multm_qsp89 & multm_qcp88;
  assign multm_compress_add3b_maj3b_wx89 = multm_qsp90 & multm_qcp89;
  assign multm_compress_add3b_maj3b_wx90 = multm_qsp91 & multm_qcp90;
  assign multm_compress_add3b_maj3b_wx91 = multm_qsp92 & multm_qcp91;
  assign multm_compress_add3b_maj3b_wx92 = multm_qsp93 & multm_qcp92;
  assign multm_compress_add3b_maj3b_wx93 = multm_qsp94 & multm_qcp93;
  assign multm_compress_add3b_maj3b_wx94 = multm_qsp95 & multm_qcp94;
  assign multm_compress_add3b_maj3b_wx95 = multm_qsp96 & multm_qcp95;
  assign multm_compress_add3b_maj3b_wx96 = multm_qsp97 & multm_qcp96;
  assign multm_compress_add3b_maj3b_wx97 = multm_qsp98 & multm_qcp97;
  assign multm_compress_add3b_maj3b_wx98 = multm_qsp99 & multm_qcp98;
  assign multm_compress_add3b_maj3b_wx99 = multm_qsp100 & multm_qcp99;
  assign multm_compress_add3b_maj3b_wx100 = multm_qsp101 & multm_qcp100;
  assign multm_compress_add3b_maj3b_wx103 = multm_qsp104 & multm_qcp103;
  assign multm_compress_add3b_maj3b_wx104 = multm_qsp105 & multm_qcp104;
  assign multm_compress_add3b_maj3b_wx106 = multm_qsp107 & multm_qcp106;
  assign multm_compress_add3b_maj3b_wx107 = multm_qsp108 & multm_qcp107;
  assign multm_compress_add3b_maj3b_wx111 = multm_qsp112 & multm_qcp111;
  assign multm_compress_add3b_maj3b_wx112 = multm_qsp113 & multm_qcp112;
  assign multm_compress_add3b_maj3b_wx113 = multm_qsp114 & multm_qcp113;
  assign multm_compress_add3b_maj3b_wx114 = multm_qsp115 & multm_qcp114;
  assign multm_compress_add3b_maj3b_wx115 = multm_qsp116 & multm_qcp115;
  assign multm_compress_add3b_maj3b_wx116 = multm_qsp117 & multm_qcp116;
  assign multm_compress_add3b_maj3b_wx117 = multm_qsp118 & multm_qcp117;
  assign multm_compress_add3b_maj3b_wx118 = multm_qsp119 & multm_qcp118;
  assign multm_compress_add3b_maj3b_wx124 = multm_qsp125 & multm_qcp124;
  assign multm_compress_add3b_maj3b_wx125 = multm_qsp126 & multm_qcp125;
  assign multm_compress_add3b_maj3b_wx126 = multm_qsp127 & multm_qcp126;
  assign multm_compress_add3b_maj3b_wx127 = multm_qsp128 & multm_qcp127;
  assign multm_compress_add3b_maj3b_wx128 = multm_qsp129 & multm_qcp128;
  assign multm_compress_add3b_maj3b_wx129 = multm_qsp130 & multm_qcp129;
  assign multm_compress_add3b_maj3b_wx130 = multm_qsp131 & multm_qcp130;
  assign multm_compress_add3b_maj3b_wx131 = multm_qsp132 & multm_qcp131;
  assign multm_compress_add3b_maj3b_wx132 = multm_qsp133 & multm_qcp132;
  assign multm_compress_add3b_maj3b_wx133 = multm_qsp134 & multm_qcp133;
  assign multm_compress_add3b_maj3b_wx134 = multm_qsp135 & multm_qcp134;
  assign multm_compress_add3b_maj3b_wx135 = multm_qsp136 & multm_qcp135;
  assign multm_compress_add3b_maj3b_wx136 = multm_qsp137 & multm_qcp136;
  assign multm_compress_add3b_maj3b_wx137 = multm_qsp138 & multm_qcp137;
  assign multm_compress_add3b_maj3b_wx138 = multm_qsp139 & multm_qcp138;
  assign multm_compress_add3b_maj3b_wx139 = multm_qsp140 & multm_qcp139;
  assign multm_compress_add3b_maj3b_wx140 = multm_qsp141 & multm_qcp140;
  assign multm_compress_add3b_maj3b_wx141 = multm_qsp142 & multm_qcp141;
  assign multm_compress_add3b_maj3b_wx145 = multm_qsp146 & multm_qcp145;
  assign multm_compress_add3b_maj3b_wx146 = multm_qsp147 & multm_qcp146;
  assign multm_compress_add3b_maj3b_wx147 = multm_qsp148 & multm_qcp147;
  assign multm_compress_add3b_maj3b_wx148 = multm_qsp149 & multm_qcp148;
  assign multm_compress_add3b_maj3b_wx149 = multm_qsp150 & multm_qcp149;
  assign multm_compress_add3b_maj3b_wx150 = multm_qsp151 & multm_qcp150;
  assign multm_compress_add3b_maj3b_wx151 = multm_qsp152 & multm_qcp151;
  assign multm_compress_add3b_maj3b_wx154 = multm_qsp155 & multm_qcp154;
  assign multm_compress_add3b_maj3b_wx155 = multm_qsp156 & multm_qcp155;
  assign multm_compress_add3b_maj3b_wx161 = multm_qsp162 & multm_qcp161;
  assign multm_compress_add3b_maj3b_wx162 = multm_qsp163 & multm_qcp162;
  assign multm_compress_add3b_maj3b_wx163 = multm_qsp164 & multm_qcp163;
  assign multm_compress_add3b_maj3b_wx164 = multm_qsp165 & multm_qcp164;
  assign multm_compress_add3b_maj3b_wx165 = multm_qsp166 & multm_qcp165;
  assign multm_compress_add3b_maj3b_wx166 = multm_qsp167 & multm_qcp166;
  assign multm_compress_add3b_maj3b_wx167 = multm_qsp168 & multm_qcp167;
  assign multm_compress_add3b_maj3b_wx168 = multm_qsp169 & multm_qcp168;
  assign multm_compress_add3b_maj3b_wx169 = multm_qsp170 & multm_qcp169;
  assign multm_compress_add3b_maj3b_wx170 = multm_qsp171 & multm_qcp170;
  assign multm_compress_add3b_maj3b_wx171 = multm_qsp172 & multm_qcp171;
  assign multm_compress_add3b_maj3b_wx172 = multm_qsp173 & multm_qcp172;
  assign multm_compress_add3b_maj3b_wx176 = multm_qsp177 & multm_qcp176;
  assign multm_compress_add3b_maj3b_wx177 = multm_qsp178 & multm_qcp177;
  assign multm_compress_add3b_maj3b_wx178 = multm_qsp179 & multm_qcp178;
  assign multm_compress_add3b_maj3b_wx179 = multm_qsp180 & multm_qcp179;
  assign multm_compress_add3b_maj3b_wx180 = multm_qsp181 & multm_qcp180;
  assign multm_compress_add3b_maj3b_wx181 = multm_qsp182 & multm_qcp181;
  assign multm_compress_add3b_maj3b_wx182 = multm_qsp183 & multm_qcp182;
  assign multm_compress_add3b_maj3b_wy0 = multm_qsp1 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_wy2 = multm_qsp3 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy3 = multm_qsp4 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy4 = multm_qsp5 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy5 = multm_qsp6 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy8 = multm_qsp9 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy9 = multm_qsp10 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy10 = multm_qsp11 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy11 = multm_qsp12 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy12 = multm_qsp13 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy13 = multm_qsp14 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy14 = multm_qsp15 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy15 = multm_qsp16 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy16 = multm_qsp17 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy17 = multm_qsp18 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy18 = multm_qsp19 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy19 = multm_qsp20 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy20 = multm_qsp21 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy21 = multm_qsp22 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy22 = multm_qsp23 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy23 = multm_qsp24 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy25 = multm_qsp26 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy26 = multm_qsp27 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy27 = multm_qsp28 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy28 = multm_qsp29 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy29 = multm_qsp30 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy30 = multm_qsp31 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy31 = multm_qsp32 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy32 = multm_qsp33 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy33 = multm_qsp34 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy34 = multm_qsp35 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy35 = multm_qsp36 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy36 = multm_qsp37 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy37 = multm_qsp38 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy38 = multm_qsp39 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy39 = multm_qsp40 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy40 = multm_qsp41 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy41 = multm_qsp42 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy44 = multm_qsp45 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy45 = multm_qsp46 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy46 = multm_qsp47 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy47 = multm_qsp48 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy48 = multm_qsp49 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy49 = multm_qsp50 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy50 = multm_qsp51 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy51 = multm_qsp52 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy52 = multm_qsp53 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy56 = multm_qsp57 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy57 = multm_qsp58 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_wy58 = multm_qsp59 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy59 = multm_qsp60 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy60 = multm_qsp61 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy61 = multm_qsp62 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy62 = multm_qsp63 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy63 = multm_qsp64 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy64 = multm_qsp65 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy65 = multm_qsp66 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy66 = multm_qsp67 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy67 = multm_qsp68 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy68 = multm_qsp69 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy69 = multm_qsp70 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy70 = multm_qsp71 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy71 = multm_qsp72 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_wy72 = multm_qsp73 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy73 = multm_qsp74 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_wy75 = multm_qsp76 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy76 = multm_qsp77 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy77 = multm_qsp78 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy78 = multm_qsp79 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy79 = multm_qsp80 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy80 = multm_qsp81 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy81 = multm_qsp82 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy82 = multm_qsp83 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_wy83 = multm_qsp84 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy84 = multm_qsp85 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy85 = multm_qsp86 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy86 = multm_qsp87 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy87 = multm_qsp88 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy88 = multm_qsp89 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy89 = multm_qsp90 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy90 = multm_qsp91 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy91 = multm_qsp92 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy92 = multm_qsp93 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy93 = multm_qsp94 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy94 = multm_qsp95 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy95 = multm_qsp96 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy96 = multm_qsp97 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy97 = multm_qsp98 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy98 = multm_qsp99 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy99 = multm_qsp100 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy100 = multm_qsp101 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy103 = multm_qsp104 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy104 = multm_qsp105 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_wy106 = multm_qsp107 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy107 = multm_qsp108 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_wy111 = multm_qsp112 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy112 = multm_qsp113 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_wy113 = multm_qsp114 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy114 = multm_qsp115 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_wy115 = multm_qsp116 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy116 = multm_qsp117 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy117 = multm_qsp118 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy118 = multm_qsp119 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy124 = multm_qsp125 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy125 = multm_qsp126 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy126 = multm_qsp127 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy127 = multm_qsp128 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy128 = multm_qsp129 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy129 = multm_qsp130 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy130 = multm_qsp131 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy131 = multm_qsp132 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy132 = multm_qsp133 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy133 = multm_qsp134 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy134 = multm_qsp135 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy135 = multm_qsp136 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy136 = multm_qsp137 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy137 = multm_qsp138 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy138 = multm_qsp139 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy139 = multm_qsp140 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy140 = multm_qsp141 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy141 = multm_qsp142 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy145 = multm_qsp146 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy146 = multm_qsp147 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy147 = multm_qsp148 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy148 = multm_qsp149 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy149 = multm_qsp150 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy150 = multm_qsp151 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy151 = multm_qsp152 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy154 = multm_qsp155 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy155 = multm_qsp156 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_wy161 = multm_qsp162 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy162 = multm_qsp163 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_wy163 = multm_qsp164 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy164 = multm_qsp165 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy165 = multm_qsp166 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy166 = multm_qsp167 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy167 = multm_qsp168 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy168 = multm_qsp169 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy169 = multm_qsp170 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy170 = multm_qsp171 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy171 = multm_qsp172 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy172 = multm_qsp173 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_wy176 = multm_qsp177 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_wy177 = multm_qsp178 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_wy178 = multm_qsp179 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_wy179 = multm_qsp180 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy180 = multm_qsp181 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_wy181 = multm_qsp182 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_wy182 = multm_qsp183 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy0 = multm_qcp0 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_xy2 = multm_qcp2 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy3 = multm_qcp3 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy4 = multm_qcp4 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy5 = multm_qcp5 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy8 = multm_qcp8 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy9 = multm_qcp9 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy10 = multm_qcp10 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy11 = multm_qcp11 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy12 = multm_qcp12 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy13 = multm_qcp13 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy14 = multm_qcp14 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy15 = multm_qcp15 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy16 = multm_qcp16 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy17 = multm_qcp17 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy18 = multm_qcp18 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy19 = multm_qcp19 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy20 = multm_qcp20 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy21 = multm_qcp21 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy22 = multm_qcp22 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy23 = multm_qcp23 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy25 = multm_qcp25 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy26 = multm_qcp26 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy27 = multm_qcp27 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy28 = multm_qcp28 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy29 = multm_qcp29 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy30 = multm_qcp30 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy31 = multm_qcp31 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy32 = multm_qcp32 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy33 = multm_qcp33 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy34 = multm_qcp34 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy35 = multm_qcp35 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy36 = multm_qcp36 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy37 = multm_qcp37 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy38 = multm_qcp38 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy39 = multm_qcp39 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy40 = multm_qcp40 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy41 = multm_qcp41 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy44 = multm_qcp44 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy45 = multm_qcp45 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy46 = multm_qcp46 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy47 = multm_qcp47 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy48 = multm_qcp48 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy49 = multm_qcp49 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy50 = multm_qcp50 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy51 = multm_qcp51 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy52 = multm_qcp52 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy56 = multm_qcp56 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy57 = multm_qcp57 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_xy58 = multm_qcp58 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy59 = multm_qcp59 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy60 = multm_qcp60 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy61 = multm_qcp61 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy62 = multm_qcp62 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy63 = multm_qcp63 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy64 = multm_qcp64 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy65 = multm_qcp65 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy66 = multm_qcp66 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy67 = multm_qcp67 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy68 = multm_qcp68 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy69 = multm_qcp69 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy70 = multm_qcp70 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy71 = multm_qcp71 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_xy72 = multm_qcp72 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy73 = multm_qcp73 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_xy75 = multm_qcp75 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy76 = multm_qcp76 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy77 = multm_qcp77 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy78 = multm_qcp78 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy79 = multm_qcp79 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy80 = multm_qcp80 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy81 = multm_qcp81 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy82 = multm_qcp82 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_xy83 = multm_qcp83 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy84 = multm_qcp84 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy85 = multm_qcp85 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy86 = multm_qcp86 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy87 = multm_qcp87 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy88 = multm_qcp88 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy89 = multm_qcp89 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy90 = multm_qcp90 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy91 = multm_qcp91 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy92 = multm_qcp92 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy93 = multm_qcp93 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy94 = multm_qcp94 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy95 = multm_qcp95 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy96 = multm_qcp96 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy97 = multm_qcp97 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy98 = multm_qcp98 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy99 = multm_qcp99 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy100 = multm_qcp100 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy103 = multm_qcp103 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy104 = multm_qcp104 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_xy106 = multm_qcp106 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy107 = multm_qcp107 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_xy111 = multm_qcp111 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy112 = multm_qcp112 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_xy113 = multm_qcp113 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy114 = multm_qcp114 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_xy115 = multm_qcp115 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy116 = multm_qcp116 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy117 = multm_qcp117 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy118 = multm_qcp118 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy124 = multm_qcp124 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy125 = multm_qcp125 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy126 = multm_qcp126 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy127 = multm_qcp127 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy128 = multm_qcp128 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy129 = multm_qcp129 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy130 = multm_qcp130 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy131 = multm_qcp131 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy132 = multm_qcp132 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy133 = multm_qcp133 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy134 = multm_qcp134 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy135 = multm_qcp135 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy136 = multm_qcp136 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy137 = multm_qcp137 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy138 = multm_qcp138 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy139 = multm_qcp139 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy140 = multm_qcp140 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy141 = multm_qcp141 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy145 = multm_qcp145 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy146 = multm_qcp146 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy147 = multm_qcp147 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy148 = multm_qcp148 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy149 = multm_qcp149 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy150 = multm_qcp150 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy151 = multm_qcp151 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy154 = multm_qcp154 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy155 = multm_qcp155 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_xy161 = multm_qcp161 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy162 = multm_qcp162 & multm_compress_ncd;
  assign multm_compress_add3b_maj3b_xy163 = multm_qcp163 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy164 = multm_qcp164 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy165 = multm_qcp165 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy166 = multm_qcp166 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy167 = multm_qcp167 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy168 = multm_qcp168 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy169 = multm_qcp169 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy170 = multm_qcp170 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy171 = multm_qcp171 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy172 = multm_qcp172 & multm_compress_rn6;
  assign multm_compress_add3b_maj3b_xy176 = multm_qcp176 & multm_compress_nsd;
  assign multm_compress_add3b_maj3b_xy177 = multm_qcp177 & multm_compress_rn4;
  assign multm_compress_add3b_maj3b_xy178 = multm_qcp178 & multm_compress_rn15;
  assign multm_compress_add3b_maj3b_xy179 = multm_qcp179 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy180 = multm_qcp180 & multm_compress_rn20;
  assign multm_compress_add3b_maj3b_xy181 = multm_qcp181 & multm_compress_rn5;
  assign multm_compress_add3b_maj3b_xy182 = multm_qcp182 & multm_compress_rn6;
  assign multm_compress_add3b_xor3b_wx0 = multm_qsp1 ^ multm_qcp0;
  assign multm_compress_add3b_xor3b_wx2 = multm_qsp3 ^ multm_qcp2;
  assign multm_compress_add3b_xor3b_wx3 = multm_qsp4 ^ multm_qcp3;
  assign multm_compress_add3b_xor3b_wx4 = multm_qsp5 ^ multm_qcp4;
  assign multm_compress_add3b_xor3b_wx5 = multm_qsp6 ^ multm_qcp5;
  assign multm_compress_add3b_xor3b_wx8 = multm_qsp9 ^ multm_qcp8;
  assign multm_compress_add3b_xor3b_wx9 = multm_qsp10 ^ multm_qcp9;
  assign multm_compress_add3b_xor3b_wx10 = multm_qsp11 ^ multm_qcp10;
  assign multm_compress_add3b_xor3b_wx11 = multm_qsp12 ^ multm_qcp11;
  assign multm_compress_add3b_xor3b_wx12 = multm_qsp13 ^ multm_qcp12;
  assign multm_compress_add3b_xor3b_wx13 = multm_qsp14 ^ multm_qcp13;
  assign multm_compress_add3b_xor3b_wx14 = multm_qsp15 ^ multm_qcp14;
  assign multm_compress_add3b_xor3b_wx15 = multm_qsp16 ^ multm_qcp15;
  assign multm_compress_add3b_xor3b_wx16 = multm_qsp17 ^ multm_qcp16;
  assign multm_compress_add3b_xor3b_wx17 = multm_qsp18 ^ multm_qcp17;
  assign multm_compress_add3b_xor3b_wx18 = multm_qsp19 ^ multm_qcp18;
  assign multm_compress_add3b_xor3b_wx19 = multm_qsp20 ^ multm_qcp19;
  assign multm_compress_add3b_xor3b_wx20 = multm_qsp21 ^ multm_qcp20;
  assign multm_compress_add3b_xor3b_wx21 = multm_qsp22 ^ multm_qcp21;
  assign multm_compress_add3b_xor3b_wx22 = multm_qsp23 ^ multm_qcp22;
  assign multm_compress_add3b_xor3b_wx23 = multm_qsp24 ^ multm_qcp23;
  assign multm_compress_add3b_xor3b_wx25 = multm_qsp26 ^ multm_qcp25;
  assign multm_compress_add3b_xor3b_wx26 = multm_qsp27 ^ multm_qcp26;
  assign multm_compress_add3b_xor3b_wx27 = multm_qsp28 ^ multm_qcp27;
  assign multm_compress_add3b_xor3b_wx28 = multm_qsp29 ^ multm_qcp28;
  assign multm_compress_add3b_xor3b_wx29 = multm_qsp30 ^ multm_qcp29;
  assign multm_compress_add3b_xor3b_wx30 = multm_qsp31 ^ multm_qcp30;
  assign multm_compress_add3b_xor3b_wx31 = multm_qsp32 ^ multm_qcp31;
  assign multm_compress_add3b_xor3b_wx32 = multm_qsp33 ^ multm_qcp32;
  assign multm_compress_add3b_xor3b_wx33 = multm_qsp34 ^ multm_qcp33;
  assign multm_compress_add3b_xor3b_wx34 = multm_qsp35 ^ multm_qcp34;
  assign multm_compress_add3b_xor3b_wx35 = multm_qsp36 ^ multm_qcp35;
  assign multm_compress_add3b_xor3b_wx36 = multm_qsp37 ^ multm_qcp36;
  assign multm_compress_add3b_xor3b_wx37 = multm_qsp38 ^ multm_qcp37;
  assign multm_compress_add3b_xor3b_wx38 = multm_qsp39 ^ multm_qcp38;
  assign multm_compress_add3b_xor3b_wx39 = multm_qsp40 ^ multm_qcp39;
  assign multm_compress_add3b_xor3b_wx40 = multm_qsp41 ^ multm_qcp40;
  assign multm_compress_add3b_xor3b_wx41 = multm_qsp42 ^ multm_qcp41;
  assign multm_compress_add3b_xor3b_wx44 = multm_qsp45 ^ multm_qcp44;
  assign multm_compress_add3b_xor3b_wx45 = multm_qsp46 ^ multm_qcp45;
  assign multm_compress_add3b_xor3b_wx46 = multm_qsp47 ^ multm_qcp46;
  assign multm_compress_add3b_xor3b_wx47 = multm_qsp48 ^ multm_qcp47;
  assign multm_compress_add3b_xor3b_wx48 = multm_qsp49 ^ multm_qcp48;
  assign multm_compress_add3b_xor3b_wx49 = multm_qsp50 ^ multm_qcp49;
  assign multm_compress_add3b_xor3b_wx50 = multm_qsp51 ^ multm_qcp50;
  assign multm_compress_add3b_xor3b_wx51 = multm_qsp52 ^ multm_qcp51;
  assign multm_compress_add3b_xor3b_wx52 = multm_qsp53 ^ multm_qcp52;
  assign multm_compress_add3b_xor3b_wx56 = multm_qsp57 ^ multm_qcp56;
  assign multm_compress_add3b_xor3b_wx57 = multm_qsp58 ^ multm_qcp57;
  assign multm_compress_add3b_xor3b_wx58 = multm_qsp59 ^ multm_qcp58;
  assign multm_compress_add3b_xor3b_wx59 = multm_qsp60 ^ multm_qcp59;
  assign multm_compress_add3b_xor3b_wx60 = multm_qsp61 ^ multm_qcp60;
  assign multm_compress_add3b_xor3b_wx61 = multm_qsp62 ^ multm_qcp61;
  assign multm_compress_add3b_xor3b_wx62 = multm_qsp63 ^ multm_qcp62;
  assign multm_compress_add3b_xor3b_wx63 = multm_qsp64 ^ multm_qcp63;
  assign multm_compress_add3b_xor3b_wx64 = multm_qsp65 ^ multm_qcp64;
  assign multm_compress_add3b_xor3b_wx65 = multm_qsp66 ^ multm_qcp65;
  assign multm_compress_add3b_xor3b_wx66 = multm_qsp67 ^ multm_qcp66;
  assign multm_compress_add3b_xor3b_wx67 = multm_qsp68 ^ multm_qcp67;
  assign multm_compress_add3b_xor3b_wx68 = multm_qsp69 ^ multm_qcp68;
  assign multm_compress_add3b_xor3b_wx69 = multm_qsp70 ^ multm_qcp69;
  assign multm_compress_add3b_xor3b_wx70 = multm_qsp71 ^ multm_qcp70;
  assign multm_compress_add3b_xor3b_wx71 = multm_qsp72 ^ multm_qcp71;
  assign multm_compress_add3b_xor3b_wx72 = multm_qsp73 ^ multm_qcp72;
  assign multm_compress_add3b_xor3b_wx73 = multm_qsp74 ^ multm_qcp73;
  assign multm_compress_add3b_xor3b_wx75 = multm_qsp76 ^ multm_qcp75;
  assign multm_compress_add3b_xor3b_wx76 = multm_qsp77 ^ multm_qcp76;
  assign multm_compress_add3b_xor3b_wx77 = multm_qsp78 ^ multm_qcp77;
  assign multm_compress_add3b_xor3b_wx78 = multm_qsp79 ^ multm_qcp78;
  assign multm_compress_add3b_xor3b_wx79 = multm_qsp80 ^ multm_qcp79;
  assign multm_compress_add3b_xor3b_wx80 = multm_qsp81 ^ multm_qcp80;
  assign multm_compress_add3b_xor3b_wx81 = multm_qsp82 ^ multm_qcp81;
  assign multm_compress_add3b_xor3b_wx82 = multm_qsp83 ^ multm_qcp82;
  assign multm_compress_add3b_xor3b_wx83 = multm_qsp84 ^ multm_qcp83;
  assign multm_compress_add3b_xor3b_wx84 = multm_qsp85 ^ multm_qcp84;
  assign multm_compress_add3b_xor3b_wx85 = multm_qsp86 ^ multm_qcp85;
  assign multm_compress_add3b_xor3b_wx86 = multm_qsp87 ^ multm_qcp86;
  assign multm_compress_add3b_xor3b_wx87 = multm_qsp88 ^ multm_qcp87;
  assign multm_compress_add3b_xor3b_wx88 = multm_qsp89 ^ multm_qcp88;
  assign multm_compress_add3b_xor3b_wx89 = multm_qsp90 ^ multm_qcp89;
  assign multm_compress_add3b_xor3b_wx90 = multm_qsp91 ^ multm_qcp90;
  assign multm_compress_add3b_xor3b_wx91 = multm_qsp92 ^ multm_qcp91;
  assign multm_compress_add3b_xor3b_wx92 = multm_qsp93 ^ multm_qcp92;
  assign multm_compress_add3b_xor3b_wx93 = multm_qsp94 ^ multm_qcp93;
  assign multm_compress_add3b_xor3b_wx94 = multm_qsp95 ^ multm_qcp94;
  assign multm_compress_add3b_xor3b_wx95 = multm_qsp96 ^ multm_qcp95;
  assign multm_compress_add3b_xor3b_wx96 = multm_qsp97 ^ multm_qcp96;
  assign multm_compress_add3b_xor3b_wx97 = multm_qsp98 ^ multm_qcp97;
  assign multm_compress_add3b_xor3b_wx98 = multm_qsp99 ^ multm_qcp98;
  assign multm_compress_add3b_xor3b_wx99 = multm_qsp100 ^ multm_qcp99;
  assign multm_compress_add3b_xor3b_wx100 = multm_qsp101 ^ multm_qcp100;
  assign multm_compress_add3b_xor3b_wx103 = multm_qsp104 ^ multm_qcp103;
  assign multm_compress_add3b_xor3b_wx104 = multm_qsp105 ^ multm_qcp104;
  assign multm_compress_add3b_xor3b_wx106 = multm_qsp107 ^ multm_qcp106;
  assign multm_compress_add3b_xor3b_wx107 = multm_qsp108 ^ multm_qcp107;
  assign multm_compress_add3b_xor3b_wx111 = multm_qsp112 ^ multm_qcp111;
  assign multm_compress_add3b_xor3b_wx112 = multm_qsp113 ^ multm_qcp112;
  assign multm_compress_add3b_xor3b_wx113 = multm_qsp114 ^ multm_qcp113;
  assign multm_compress_add3b_xor3b_wx114 = multm_qsp115 ^ multm_qcp114;
  assign multm_compress_add3b_xor3b_wx115 = multm_qsp116 ^ multm_qcp115;
  assign multm_compress_add3b_xor3b_wx116 = multm_qsp117 ^ multm_qcp116;
  assign multm_compress_add3b_xor3b_wx117 = multm_qsp118 ^ multm_qcp117;
  assign multm_compress_add3b_xor3b_wx118 = multm_qsp119 ^ multm_qcp118;
  assign multm_compress_add3b_xor3b_wx124 = multm_qsp125 ^ multm_qcp124;
  assign multm_compress_add3b_xor3b_wx125 = multm_qsp126 ^ multm_qcp125;
  assign multm_compress_add3b_xor3b_wx126 = multm_qsp127 ^ multm_qcp126;
  assign multm_compress_add3b_xor3b_wx127 = multm_qsp128 ^ multm_qcp127;
  assign multm_compress_add3b_xor3b_wx128 = multm_qsp129 ^ multm_qcp128;
  assign multm_compress_add3b_xor3b_wx129 = multm_qsp130 ^ multm_qcp129;
  assign multm_compress_add3b_xor3b_wx130 = multm_qsp131 ^ multm_qcp130;
  assign multm_compress_add3b_xor3b_wx131 = multm_qsp132 ^ multm_qcp131;
  assign multm_compress_add3b_xor3b_wx132 = multm_qsp133 ^ multm_qcp132;
  assign multm_compress_add3b_xor3b_wx133 = multm_qsp134 ^ multm_qcp133;
  assign multm_compress_add3b_xor3b_wx134 = multm_qsp135 ^ multm_qcp134;
  assign multm_compress_add3b_xor3b_wx135 = multm_qsp136 ^ multm_qcp135;
  assign multm_compress_add3b_xor3b_wx136 = multm_qsp137 ^ multm_qcp136;
  assign multm_compress_add3b_xor3b_wx137 = multm_qsp138 ^ multm_qcp137;
  assign multm_compress_add3b_xor3b_wx138 = multm_qsp139 ^ multm_qcp138;
  assign multm_compress_add3b_xor3b_wx139 = multm_qsp140 ^ multm_qcp139;
  assign multm_compress_add3b_xor3b_wx140 = multm_qsp141 ^ multm_qcp140;
  assign multm_compress_add3b_xor3b_wx141 = multm_qsp142 ^ multm_qcp141;
  assign multm_compress_add3b_xor3b_wx145 = multm_qsp146 ^ multm_qcp145;
  assign multm_compress_add3b_xor3b_wx146 = multm_qsp147 ^ multm_qcp146;
  assign multm_compress_add3b_xor3b_wx147 = multm_qsp148 ^ multm_qcp147;
  assign multm_compress_add3b_xor3b_wx148 = multm_qsp149 ^ multm_qcp148;
  assign multm_compress_add3b_xor3b_wx149 = multm_qsp150 ^ multm_qcp149;
  assign multm_compress_add3b_xor3b_wx150 = multm_qsp151 ^ multm_qcp150;
  assign multm_compress_add3b_xor3b_wx151 = multm_qsp152 ^ multm_qcp151;
  assign multm_compress_add3b_xor3b_wx154 = multm_qsp155 ^ multm_qcp154;
  assign multm_compress_add3b_xor3b_wx155 = multm_qsp156 ^ multm_qcp155;
  assign multm_compress_add3b_xor3b_wx161 = multm_qsp162 ^ multm_qcp161;
  assign multm_compress_add3b_xor3b_wx162 = multm_qsp163 ^ multm_qcp162;
  assign multm_compress_add3b_xor3b_wx163 = multm_qsp164 ^ multm_qcp163;
  assign multm_compress_add3b_xor3b_wx164 = multm_qsp165 ^ multm_qcp164;
  assign multm_compress_add3b_xor3b_wx165 = multm_qsp166 ^ multm_qcp165;
  assign multm_compress_add3b_xor3b_wx166 = multm_qsp167 ^ multm_qcp166;
  assign multm_compress_add3b_xor3b_wx167 = multm_qsp168 ^ multm_qcp167;
  assign multm_compress_add3b_xor3b_wx168 = multm_qsp169 ^ multm_qcp168;
  assign multm_compress_add3b_xor3b_wx169 = multm_qsp170 ^ multm_qcp169;
  assign multm_compress_add3b_xor3b_wx170 = multm_qsp171 ^ multm_qcp170;
  assign multm_compress_add3b_xor3b_wx171 = multm_qsp172 ^ multm_qcp171;
  assign multm_compress_add3b_xor3b_wx172 = multm_qsp173 ^ multm_qcp172;
  assign multm_compress_add3b_xor3b_wx176 = multm_qsp177 ^ multm_qcp176;
  assign multm_compress_add3b_xor3b_wx177 = multm_qsp178 ^ multm_qcp177;
  assign multm_compress_add3b_xor3b_wx178 = multm_qsp179 ^ multm_qcp178;
  assign multm_compress_add3b_xor3b_wx179 = multm_qsp180 ^ multm_qcp179;
  assign multm_compress_add3b_xor3b_wx180 = multm_qsp181 ^ multm_qcp180;
  assign multm_compress_add3b_xor3b_wx181 = multm_qsp182 ^ multm_qcp181;
  assign multm_compress_add3b_xor3b_wx182 = multm_qsp183 ^ multm_qcp182;
  assign multm_compress_nc = multm_compress_nct | multm_qcp184;
  assign multm_compress_nct = multm_qsp184 & multm_qcp183;
  assign multm_compress_ns = multm_qsp184 ^ multm_qcp183;
  assign multm_compress_rn4 = multm_compress_ncd ? multm_compress_rnh4 : multm_compress_nsd;
  assign multm_compress_rn5 = multm_compress_ncd & multm_compress_rnh4;
  assign multm_compress_rn6 = multm_compress_ncd & multm_compress_nsd;
  assign multm_compress_rn15 = multm_compress_ncd | multm_compress_nsd;
  assign multm_compress_rn20 = xn6 & multm_compress_nsd;
  assign multm_compress_rnh4 = ~multm_compress_nsd;
  assign multm_ctrp_ctr_cq0 = ~multm_ctrp_ctr_cp0;
  assign multm_ctrp_ctr_cq1 = multm_ctrp_ctr_sp0 & multm_ctrp_ctr_cp0;
  assign multm_ctrp_ctr_cq2 = multm_ctrp_ctr_sp1 & multm_ctrp_ctr_cp1;
  assign multm_ctrp_ctr_cq3 = multm_ctrp_ctr_sp2 & multm_ctrp_ctr_cp2;
  assign multm_ctrp_ctr_cq4 = multm_ctrp_ctr_sp3 & multm_ctrp_ctr_cp3;
  assign multm_ctrp_ctr_cq5 = multm_ctrp_ctr_sp4 & multm_ctrp_ctr_cp4;
  assign multm_ctrp_ctr_cq6 = multm_ctrp_ctr_sp5 & multm_ctrp_ctr_cp5;
  assign multm_ctrp_ctr_cq7 = multm_ctrp_ctr_sp6 & multm_ctrp_ctr_cp6;
  assign multm_ctrp_ctr_cr0 = sadd | multm_ctrp_ctr_cq0;
  assign multm_ctrp_ctr_cr1 = xn4 & multm_ctrp_ctr_cq1;
  assign multm_ctrp_ctr_cr2 = xn4 & multm_ctrp_ctr_cq2;
  assign multm_ctrp_ctr_cr3 = xn4 & multm_ctrp_ctr_cq3;
  assign multm_ctrp_ctr_cr4 = xn4 & multm_ctrp_ctr_cq4;
  assign multm_ctrp_ctr_cr5 = xn4 & multm_ctrp_ctr_cq5;
  assign multm_ctrp_ctr_cr6 = xn4 & multm_ctrp_ctr_cq6;
  assign multm_ctrp_ctr_cr7 = xn4 & multm_ctrp_ctr_cq7;
  assign multm_ctrp_ctr_dq = multm_ctrp_ctr_dp | multm_ctrp_ctr_cp7;
  assign multm_ctrp_ctr_sq0 = multm_ctrp_ctr_sp0 ^ multm_ctrp_ctr_cp0;
  assign multm_ctrp_ctr_sq1 = multm_ctrp_ctr_sp1 ^ multm_ctrp_ctr_cp1;
  assign multm_ctrp_ctr_sq2 = multm_ctrp_ctr_sp2 ^ multm_ctrp_ctr_cp2;
  assign multm_ctrp_ctr_sq3 = multm_ctrp_ctr_sp3 ^ multm_ctrp_ctr_cp3;
  assign multm_ctrp_ctr_sq4 = multm_ctrp_ctr_sp4 ^ multm_ctrp_ctr_cp4;
  assign multm_ctrp_ctr_sq5 = multm_ctrp_ctr_sp5 ^ multm_ctrp_ctr_cp5;
  assign multm_ctrp_ctr_sq6 = multm_ctrp_ctr_sp6 ^ multm_ctrp_ctr_cp6;
  assign multm_ctrp_ctr_sr0 = sadd | multm_ctrp_ctr_sq0;
  assign multm_ctrp_ctr_sr1 = xn4 & multm_ctrp_ctr_sq1;
  assign multm_ctrp_ctr_sr2 = xn4 & multm_ctrp_ctr_sq2;
  assign multm_ctrp_ctr_sr3 = xn4 & multm_ctrp_ctr_sq3;
  assign multm_ctrp_ctr_sr4 = xn4 & multm_ctrp_ctr_sq4;
  assign multm_ctrp_ctr_sr5 = sadd | multm_ctrp_ctr_sq5;
  assign multm_ctrp_ctr_sr6 = xn4 & multm_ctrp_ctr_sq6;
  assign multm_ctrp_ds = xn4 & multm_ctrp_ctr_dq;
  assign multm_ctrp_pulse_xn = ~multm_ctrp_ctr_dp;
  assign multm_pc0 = multm_reduce_add3b0_maj3b_or3b_wx0 | multm_reduce_add3b0_maj3b_xy0;
  assign multm_pc1 = multm_reduce_add3b0_maj3b_or3b_wx1 | multm_reduce_add3b0_maj3b_xy1;
  assign multm_pc2 = multm_reduce_add3b0_maj3b_or3b_wx2 | multm_reduce_add3b0_maj3b_xy2;
  assign multm_pc3 = multm_reduce_add3b0_maj3b_or3b_wx3 | multm_reduce_add3b0_maj3b_xy3;
  assign multm_pc4 = multm_reduce_add3b0_maj3b_or3b_wx4 | multm_reduce_add3b0_maj3b_xy4;
  assign multm_pc5 = multm_reduce_add3b0_maj3b_or3b_wx5 | multm_reduce_add3b0_maj3b_xy5;
  assign multm_pc6 = multm_reduce_add3b0_maj3b_or3b_wx6 | multm_reduce_add3b0_maj3b_xy6;
  assign multm_pc7 = multm_reduce_add3b0_maj3b_or3b_wx7 | multm_reduce_add3b0_maj3b_xy7;
  assign multm_pc8 = multm_reduce_add3b0_maj3b_or3b_wx8 | multm_reduce_add3b0_maj3b_xy8;
  assign multm_pc9 = multm_reduce_add3b0_maj3b_or3b_wx9 | multm_reduce_add3b0_maj3b_xy9;
  assign multm_pc11 = multm_reduce_add3b1_maj3b_or3b_wx0 | multm_reduce_add3b1_maj3b_xy0;
  assign multm_pc12 = multm_reduce_add3b1_maj3b_or3b_wx1 | multm_reduce_add3b1_maj3b_xy1;
  assign multm_pc13 = multm_reduce_add3b1_maj3b_or3b_wx2 | multm_reduce_add3b1_maj3b_xy2;
  assign multm_pc14 = multm_reduce_add3b1_maj3b_or3b_wx3 | multm_reduce_add3b1_maj3b_xy3;
  assign multm_pc15 = multm_reduce_add3b1_maj3b_or3b_wx4 | multm_reduce_add3b1_maj3b_xy4;
  assign multm_pc16 = multm_reduce_add3b1_maj3b_or3b_wx5 | multm_reduce_add3b1_maj3b_xy5;
  assign multm_pc17 = multm_reduce_add3b1_maj3b_or3b_wx6 | multm_reduce_add3b1_maj3b_xy6;
  assign multm_pc18 = multm_reduce_add3b1_maj3b_or3b_wx7 | multm_reduce_add3b1_maj3b_xy7;
  assign multm_pc19 = multm_reduce_add3b1_maj3b_or3b_wx8 | multm_reduce_add3b1_maj3b_xy8;
  assign multm_pc20 = multm_reduce_add3b1_maj3b_or3b_wx9 | multm_reduce_add3b1_maj3b_xy9;
  assign multm_pc21 = multm_reduce_add3b1_maj3b_or3b_wx10 | multm_reduce_add3b1_maj3b_xy10;
  assign multm_pc22 = multm_reduce_add3b1_maj3b_or3b_wx11 | multm_reduce_add3b1_maj3b_xy11;
  assign multm_pc23 = multm_reduce_add3b1_maj3b_or3b_wx12 | multm_reduce_add3b1_maj3b_xy12;
  assign multm_pc24 = multm_reduce_add3b1_maj3b_or3b_wx13 | multm_reduce_add3b1_maj3b_xy13;
  assign multm_pc25 = multm_reduce_add3b1_maj3b_or3b_wx14 | multm_reduce_add3b1_maj3b_xy14;
  assign multm_pc26 = multm_reduce_add3b1_maj3b_or3b_wx15 | multm_reduce_add3b1_maj3b_xy15;
  assign multm_pc27 = multm_reduce_add3b1_maj3b_or3b_wx16 | multm_reduce_add3b1_maj3b_xy16;
  assign multm_pc28 = multm_reduce_add3b1_maj3b_or3b_wx17 | multm_reduce_add3b1_maj3b_xy17;
  assign multm_pc29 = multm_reduce_add3b1_maj3b_or3b_wx18 | multm_reduce_add3b1_maj3b_xy18;
  assign multm_pc30 = multm_reduce_add3b1_maj3b_or3b_wx19 | multm_reduce_add3b1_maj3b_xy19;
  assign multm_pc31 = multm_reduce_add3b1_maj3b_or3b_wx20 | multm_reduce_add3b1_maj3b_xy20;
  assign multm_pc32 = multm_reduce_add3b1_maj3b_or3b_wx21 | multm_reduce_add3b1_maj3b_xy21;
  assign multm_pc33 = multm_reduce_add3b1_maj3b_or3b_wx22 | multm_reduce_add3b1_maj3b_xy22;
  assign multm_pc34 = multm_reduce_add3b1_maj3b_or3b_wx23 | multm_reduce_add3b1_maj3b_xy23;
  assign multm_pc35 = multm_reduce_add3b1_maj3b_or3b_wx24 | multm_reduce_add3b1_maj3b_xy24;
  assign multm_pc36 = multm_reduce_add3b1_maj3b_or3b_wx25 | multm_reduce_add3b1_maj3b_xy25;
  assign multm_pc37 = multm_reduce_add3b1_maj3b_or3b_wx26 | multm_reduce_add3b1_maj3b_xy26;
  assign multm_pc38 = multm_reduce_add3b1_maj3b_or3b_wx27 | multm_reduce_add3b1_maj3b_xy27;
  assign multm_pc39 = multm_reduce_add3b1_maj3b_or3b_wx28 | multm_reduce_add3b1_maj3b_xy28;
  assign multm_pc40 = multm_reduce_add3b1_maj3b_or3b_wx29 | multm_reduce_add3b1_maj3b_xy29;
  assign multm_pc41 = multm_reduce_add3b1_maj3b_or3b_wx30 | multm_reduce_add3b1_maj3b_xy30;
  assign multm_pc42 = multm_reduce_add3b1_maj3b_or3b_wx31 | multm_reduce_add3b1_maj3b_xy31;
  assign multm_pc43 = multm_reduce_add3b1_maj3b_or3b_wx32 | multm_reduce_add3b1_maj3b_xy32;
  assign multm_pc44 = multm_reduce_add3b1_maj3b_or3b_wx33 | multm_reduce_add3b1_maj3b_xy33;
  assign multm_pc45 = multm_reduce_add3b1_maj3b_or3b_wx34 | multm_reduce_add3b1_maj3b_xy34;
  assign multm_pc46 = multm_reduce_add3b1_maj3b_or3b_wx35 | multm_reduce_add3b1_maj3b_xy35;
  assign multm_pc47 = multm_reduce_add3b1_maj3b_or3b_wx36 | multm_reduce_add3b1_maj3b_xy36;
  assign multm_pc48 = multm_reduce_add3b1_maj3b_or3b_wx37 | multm_reduce_add3b1_maj3b_xy37;
  assign multm_pc49 = multm_reduce_add3b1_maj3b_or3b_wx38 | multm_reduce_add3b1_maj3b_xy38;
  assign multm_pc50 = multm_reduce_add3b1_maj3b_or3b_wx39 | multm_reduce_add3b1_maj3b_xy39;
  assign multm_pc51 = multm_reduce_add3b1_maj3b_or3b_wx40 | multm_reduce_add3b1_maj3b_xy40;
  assign multm_pc52 = multm_reduce_add3b1_maj3b_or3b_wx41 | multm_reduce_add3b1_maj3b_xy41;
  assign multm_pc53 = multm_reduce_add3b1_maj3b_or3b_wx42 | multm_reduce_add3b1_maj3b_xy42;
  assign multm_pc54 = multm_reduce_add3b1_maj3b_or3b_wx43 | multm_reduce_add3b1_maj3b_xy43;
  assign multm_pc55 = multm_reduce_add3b1_maj3b_or3b_wx44 | multm_reduce_add3b1_maj3b_xy44;
  assign multm_pc56 = multm_reduce_add3b1_maj3b_or3b_wx45 | multm_reduce_add3b1_maj3b_xy45;
  assign multm_pc57 = multm_reduce_add3b1_maj3b_or3b_wx46 | multm_reduce_add3b1_maj3b_xy46;
  assign multm_pc58 = multm_reduce_add3b1_maj3b_or3b_wx47 | multm_reduce_add3b1_maj3b_xy47;
  assign multm_pc59 = multm_reduce_add3b1_maj3b_or3b_wx48 | multm_reduce_add3b1_maj3b_xy48;
  assign multm_pc60 = multm_reduce_add3b1_maj3b_or3b_wx49 | multm_reduce_add3b1_maj3b_xy49;
  assign multm_pc61 = multm_reduce_add3b1_maj3b_or3b_wx50 | multm_reduce_add3b1_maj3b_xy50;
  assign multm_pc62 = multm_reduce_add3b1_maj3b_or3b_wx51 | multm_reduce_add3b1_maj3b_xy51;
  assign multm_pc63 = multm_reduce_add3b1_maj3b_or3b_wx52 | multm_reduce_add3b1_maj3b_xy52;
  assign multm_pc64 = multm_reduce_add3b1_maj3b_or3b_wx53 | multm_reduce_add3b1_maj3b_xy53;
  assign multm_pc65 = multm_reduce_add3b1_maj3b_or3b_wx54 | multm_reduce_add3b1_maj3b_xy54;
  assign multm_pc66 = multm_reduce_add3b1_maj3b_or3b_wx55 | multm_reduce_add3b1_maj3b_xy55;
  assign multm_pc67 = multm_reduce_add3b1_maj3b_or3b_wx56 | multm_reduce_add3b1_maj3b_xy56;
  assign multm_pc68 = multm_reduce_add3b1_maj3b_or3b_wx57 | multm_reduce_add3b1_maj3b_xy57;
  assign multm_pc69 = multm_reduce_add3b1_maj3b_or3b_wx58 | multm_reduce_add3b1_maj3b_xy58;
  assign multm_pc70 = multm_reduce_add3b1_maj3b_or3b_wx59 | multm_reduce_add3b1_maj3b_xy59;
  assign multm_pc71 = multm_reduce_add3b1_maj3b_or3b_wx60 | multm_reduce_add3b1_maj3b_xy60;
  assign multm_pc72 = multm_reduce_add3b1_maj3b_or3b_wx61 | multm_reduce_add3b1_maj3b_xy61;
  assign multm_pc73 = multm_reduce_add3b1_maj3b_or3b_wx62 | multm_reduce_add3b1_maj3b_xy62;
  assign multm_pc74 = multm_reduce_add3b1_maj3b_or3b_wx63 | multm_reduce_add3b1_maj3b_xy63;
  assign multm_pc75 = multm_reduce_add3b1_maj3b_or3b_wx64 | multm_reduce_add3b1_maj3b_xy64;
  assign multm_pc76 = multm_reduce_add3b1_maj3b_or3b_wx65 | multm_reduce_add3b1_maj3b_xy65;
  assign multm_pc77 = multm_reduce_add3b1_maj3b_or3b_wx66 | multm_reduce_add3b1_maj3b_xy66;
  assign multm_pc78 = multm_reduce_add3b1_maj3b_or3b_wx67 | multm_reduce_add3b1_maj3b_xy67;
  assign multm_pc79 = multm_reduce_add3b1_maj3b_or3b_wx68 | multm_reduce_add3b1_maj3b_xy68;
  assign multm_pc80 = multm_reduce_add3b1_maj3b_or3b_wx69 | multm_reduce_add3b1_maj3b_xy69;
  assign multm_pc81 = multm_reduce_add3b1_maj3b_or3b_wx70 | multm_reduce_add3b1_maj3b_xy70;
  assign multm_pc82 = multm_reduce_add3b1_maj3b_or3b_wx71 | multm_reduce_add3b1_maj3b_xy71;
  assign multm_pc83 = multm_reduce_add3b1_maj3b_or3b_wx72 | multm_reduce_add3b1_maj3b_xy72;
  assign multm_pc84 = multm_reduce_add3b1_maj3b_or3b_wx73 | multm_reduce_add3b1_maj3b_xy73;
  assign multm_pc85 = multm_reduce_add3b1_maj3b_or3b_wx74 | multm_reduce_add3b1_maj3b_xy74;
  assign multm_pc86 = multm_reduce_add3b1_maj3b_or3b_wx75 | multm_reduce_add3b1_maj3b_xy75;
  assign multm_pc87 = multm_reduce_add3b1_maj3b_or3b_wx76 | multm_reduce_add3b1_maj3b_xy76;
  assign multm_pc88 = multm_reduce_add3b1_maj3b_or3b_wx77 | multm_reduce_add3b1_maj3b_xy77;
  assign multm_pc89 = multm_reduce_add3b1_maj3b_or3b_wx78 | multm_reduce_add3b1_maj3b_xy78;
  assign multm_pc90 = multm_reduce_add3b1_maj3b_or3b_wx79 | multm_reduce_add3b1_maj3b_xy79;
  assign multm_pc91 = multm_reduce_add3b1_maj3b_or3b_wx80 | multm_reduce_add3b1_maj3b_xy80;
  assign multm_pc92 = multm_reduce_add3b1_maj3b_or3b_wx81 | multm_reduce_add3b1_maj3b_xy81;
  assign multm_pc93 = multm_reduce_add3b1_maj3b_or3b_wx82 | multm_reduce_add3b1_maj3b_xy82;
  assign multm_pc94 = multm_reduce_add3b1_maj3b_or3b_wx83 | multm_reduce_add3b1_maj3b_xy83;
  assign multm_pc95 = multm_reduce_add3b1_maj3b_or3b_wx84 | multm_reduce_add3b1_maj3b_xy84;
  assign multm_pc96 = multm_reduce_add3b1_maj3b_or3b_wx85 | multm_reduce_add3b1_maj3b_xy85;
  assign multm_pc97 = multm_reduce_add3b1_maj3b_or3b_wx86 | multm_reduce_add3b1_maj3b_xy86;
  assign multm_pc98 = multm_reduce_add3b1_maj3b_or3b_wx87 | multm_reduce_add3b1_maj3b_xy87;
  assign multm_pc99 = multm_reduce_add3b1_maj3b_or3b_wx88 | multm_reduce_add3b1_maj3b_xy88;
  assign multm_pc100 = multm_reduce_add3b1_maj3b_or3b_wx89 | multm_reduce_add3b1_maj3b_xy89;
  assign multm_pc101 = multm_reduce_add3b1_maj3b_or3b_wx90 | multm_reduce_add3b1_maj3b_xy90;
  assign multm_pc102 = multm_reduce_add3b1_maj3b_or3b_wx91 | multm_reduce_add3b1_maj3b_xy91;
  assign multm_pc103 = multm_reduce_add3b1_maj3b_or3b_wx92 | multm_reduce_add3b1_maj3b_xy92;
  assign multm_pc104 = multm_reduce_add3b1_maj3b_or3b_wx93 | multm_reduce_add3b1_maj3b_xy93;
  assign multm_pc105 = multm_reduce_add3b1_maj3b_or3b_wx94 | multm_reduce_add3b1_maj3b_xy94;
  assign multm_pc106 = multm_reduce_add3b1_maj3b_or3b_wx95 | multm_reduce_add3b1_maj3b_xy95;
  assign multm_pc107 = multm_reduce_add3b1_maj3b_or3b_wx96 | multm_reduce_add3b1_maj3b_xy96;
  assign multm_pc108 = multm_reduce_add3b1_maj3b_or3b_wx97 | multm_reduce_add3b1_maj3b_xy97;
  assign multm_pc109 = multm_reduce_add3b1_maj3b_or3b_wx98 | multm_reduce_add3b1_maj3b_xy98;
  assign multm_pc110 = multm_reduce_add3b1_maj3b_or3b_wx99 | multm_reduce_add3b1_maj3b_xy99;
  assign multm_pc111 = multm_reduce_add3b1_maj3b_or3b_wx100 | multm_reduce_add3b1_maj3b_xy100;
  assign multm_pc112 = multm_reduce_add3b1_maj3b_or3b_wx101 | multm_reduce_add3b1_maj3b_xy101;
  assign multm_pc113 = multm_reduce_add3b1_maj3b_or3b_wx102 | multm_reduce_add3b1_maj3b_xy102;
  assign multm_pc114 = multm_reduce_add3b1_maj3b_or3b_wx103 | multm_reduce_add3b1_maj3b_xy103;
  assign multm_pc115 = multm_reduce_add3b1_maj3b_or3b_wx104 | multm_reduce_add3b1_maj3b_xy104;
  assign multm_pc116 = multm_reduce_add3b1_maj3b_or3b_wx105 | multm_reduce_add3b1_maj3b_xy105;
  assign multm_pc117 = multm_reduce_add3b1_maj3b_or3b_wx106 | multm_reduce_add3b1_maj3b_xy106;
  assign multm_pc118 = multm_reduce_add3b1_maj3b_or3b_wx107 | multm_reduce_add3b1_maj3b_xy107;
  assign multm_pc119 = multm_reduce_add3b1_maj3b_or3b_wx108 | multm_reduce_add3b1_maj3b_xy108;
  assign multm_pc120 = multm_reduce_add3b1_maj3b_or3b_wx109 | multm_reduce_add3b1_maj3b_xy109;
  assign multm_pc121 = multm_reduce_add3b1_maj3b_or3b_wx110 | multm_reduce_add3b1_maj3b_xy110;
  assign multm_pc122 = multm_reduce_add3b1_maj3b_or3b_wx111 | multm_reduce_add3b1_maj3b_xy111;
  assign multm_pc123 = multm_reduce_add3b1_maj3b_or3b_wx112 | multm_reduce_add3b1_maj3b_xy112;
  assign multm_pc124 = multm_reduce_add3b1_maj3b_or3b_wx113 | multm_reduce_add3b1_maj3b_xy113;
  assign multm_pc125 = multm_reduce_add3b1_maj3b_or3b_wx114 | multm_reduce_add3b1_maj3b_xy114;
  assign multm_pc126 = multm_reduce_add3b1_maj3b_or3b_wx115 | multm_reduce_add3b1_maj3b_xy115;
  assign multm_pc127 = multm_reduce_add3b1_maj3b_or3b_wx116 | multm_reduce_add3b1_maj3b_xy116;
  assign multm_pc128 = multm_reduce_add3b1_maj3b_or3b_wx117 | multm_reduce_add3b1_maj3b_xy117;
  assign multm_pc129 = multm_reduce_add3b1_maj3b_or3b_wx118 | multm_reduce_add3b1_maj3b_xy118;
  assign multm_pc130 = multm_reduce_add3b1_maj3b_or3b_wx119 | multm_reduce_add3b1_maj3b_xy119;
  assign multm_pc131 = multm_reduce_add3b1_maj3b_or3b_wx120 | multm_reduce_add3b1_maj3b_xy120;
  assign multm_pc132 = multm_reduce_add3b1_maj3b_or3b_wx121 | multm_reduce_add3b1_maj3b_xy121;
  assign multm_pc133 = multm_reduce_add3b1_maj3b_or3b_wx122 | multm_reduce_add3b1_maj3b_xy122;
  assign multm_pc134 = multm_reduce_add3b1_maj3b_or3b_wx123 | multm_reduce_add3b1_maj3b_xy123;
  assign multm_pc135 = multm_reduce_add3b1_maj3b_or3b_wx124 | multm_reduce_add3b1_maj3b_xy124;
  assign multm_pc136 = multm_reduce_add3b1_maj3b_or3b_wx125 | multm_reduce_add3b1_maj3b_xy125;
  assign multm_pc137 = multm_reduce_add3b1_maj3b_or3b_wx126 | multm_reduce_add3b1_maj3b_xy126;
  assign multm_pc138 = multm_reduce_add3b1_maj3b_or3b_wx127 | multm_reduce_add3b1_maj3b_xy127;
  assign multm_pc139 = multm_reduce_add3b1_maj3b_or3b_wx128 | multm_reduce_add3b1_maj3b_xy128;
  assign multm_pc140 = multm_reduce_add3b1_maj3b_or3b_wx129 | multm_reduce_add3b1_maj3b_xy129;
  assign multm_pc141 = multm_reduce_add3b1_maj3b_or3b_wx130 | multm_reduce_add3b1_maj3b_xy130;
  assign multm_pc142 = multm_reduce_add3b1_maj3b_or3b_wx131 | multm_reduce_add3b1_maj3b_xy131;
  assign multm_pc143 = multm_reduce_add3b1_maj3b_or3b_wx132 | multm_reduce_add3b1_maj3b_xy132;
  assign multm_pc144 = multm_reduce_add3b1_maj3b_or3b_wx133 | multm_reduce_add3b1_maj3b_xy133;
  assign multm_pc145 = multm_reduce_add3b1_maj3b_or3b_wx134 | multm_reduce_add3b1_maj3b_xy134;
  assign multm_pc146 = multm_reduce_add3b1_maj3b_or3b_wx135 | multm_reduce_add3b1_maj3b_xy135;
  assign multm_pc147 = multm_reduce_add3b1_maj3b_or3b_wx136 | multm_reduce_add3b1_maj3b_xy136;
  assign multm_pc148 = multm_reduce_add3b1_maj3b_or3b_wx137 | multm_reduce_add3b1_maj3b_xy137;
  assign multm_pc149 = multm_reduce_add3b1_maj3b_or3b_wx138 | multm_reduce_add3b1_maj3b_xy138;
  assign multm_pc150 = multm_reduce_add3b1_maj3b_or3b_wx139 | multm_reduce_add3b1_maj3b_xy139;
  assign multm_pc151 = multm_reduce_add3b1_maj3b_or3b_wx140 | multm_reduce_add3b1_maj3b_xy140;
  assign multm_pc152 = multm_reduce_add3b1_maj3b_or3b_wx141 | multm_reduce_add3b1_maj3b_xy141;
  assign multm_pc153 = multm_reduce_add3b1_maj3b_or3b_wx142 | multm_reduce_add3b1_maj3b_xy142;
  assign multm_pc154 = multm_reduce_add3b1_maj3b_or3b_wx143 | multm_reduce_add3b1_maj3b_xy143;
  assign multm_pc155 = multm_reduce_add3b1_maj3b_or3b_wx144 | multm_reduce_add3b1_maj3b_xy144;
  assign multm_pc156 = multm_reduce_add3b1_maj3b_or3b_wx145 | multm_reduce_add3b1_maj3b_xy145;
  assign multm_pc157 = multm_reduce_add3b1_maj3b_or3b_wx146 | multm_reduce_add3b1_maj3b_xy146;
  assign multm_pc158 = multm_reduce_add3b1_maj3b_or3b_wx147 | multm_reduce_add3b1_maj3b_xy147;
  assign multm_pc159 = multm_reduce_add3b1_maj3b_or3b_wx148 | multm_reduce_add3b1_maj3b_xy148;
  assign multm_pc160 = multm_reduce_add3b1_maj3b_or3b_wx149 | multm_reduce_add3b1_maj3b_xy149;
  assign multm_pc161 = multm_reduce_add3b1_maj3b_or3b_wx150 | multm_reduce_add3b1_maj3b_xy150;
  assign multm_pc162 = multm_reduce_add3b1_maj3b_or3b_wx151 | multm_reduce_add3b1_maj3b_xy151;
  assign multm_pc163 = multm_reduce_add3b1_maj3b_or3b_wx152 | multm_reduce_add3b1_maj3b_xy152;
  assign multm_pc164 = multm_reduce_add3b1_maj3b_or3b_wx153 | multm_reduce_add3b1_maj3b_xy153;
  assign multm_pc165 = multm_reduce_add3b1_maj3b_or3b_wx154 | multm_reduce_add3b1_maj3b_xy154;
  assign multm_pc166 = multm_reduce_add3b1_maj3b_or3b_wx155 | multm_reduce_add3b1_maj3b_xy155;
  assign multm_pc167 = multm_reduce_add3b1_maj3b_or3b_wx156 | multm_reduce_add3b1_maj3b_xy156;
  assign multm_pc168 = multm_reduce_add3b1_maj3b_or3b_wx157 | multm_reduce_add3b1_maj3b_xy157;
  assign multm_pc169 = multm_reduce_add3b1_maj3b_or3b_wx158 | multm_reduce_add3b1_maj3b_xy158;
  assign multm_pc170 = multm_reduce_add3b1_maj3b_or3b_wx159 | multm_reduce_add3b1_maj3b_xy159;
  assign multm_pc171 = multm_reduce_add3b1_maj3b_or3b_wx160 | multm_reduce_add3b1_maj3b_xy160;
  assign multm_pc172 = multm_reduce_add3b1_maj3b_or3b_wx161 | multm_reduce_add3b1_maj3b_xy161;
  assign multm_pc173 = multm_reduce_add3b1_maj3b_or3b_wx162 | multm_reduce_add3b1_maj3b_xy162;
  assign multm_pc174 = multm_reduce_add3b1_maj3b_or3b_wx163 | multm_reduce_add3b1_maj3b_xy163;
  assign multm_pc175 = multm_reduce_add3b1_maj3b_or3b_wx164 | multm_reduce_add3b1_maj3b_xy164;
  assign multm_pc176 = multm_reduce_add3b1_maj3b_or3b_wx165 | multm_reduce_add3b1_maj3b_xy165;
  assign multm_pc177 = multm_reduce_add3b1_maj3b_or3b_wx166 | multm_reduce_add3b1_maj3b_xy166;
  assign multm_pc178 = multm_reduce_add3b1_maj3b_or3b_wx167 | multm_reduce_add3b1_maj3b_xy167;
  assign multm_pc179 = multm_reduce_add3b1_maj3b_or3b_wx168 | multm_reduce_add3b1_maj3b_xy168;
  assign multm_pc180 = multm_reduce_add3b1_maj3b_or3b_wx169 | multm_reduce_add3b1_maj3b_xy169;
  assign multm_pc181 = multm_reduce_add3b1_maj3b_or3b_wx170 | multm_reduce_add3b1_maj3b_xy170;
  assign multm_pc182 = multm_reduce_add3b1_maj3b_or3b_wx171 | multm_reduce_add3b1_maj3b_xy171;
  assign multm_pc183 = multm_reduce_add3b1_maj3b_or3b_wx172 | multm_reduce_add3b1_maj3b_xy172;
  assign multm_pc184 = multm_reduce_or3_wx | multm_reduce_mw;
  assign multm_ps0 = multm_reduce_add3b0_xor3b_wx0 ^ multm_reduce_sd0;
  assign multm_ps1 = multm_reduce_add3b0_xor3b_wx1 ^ multm_reduce_sd1;
  assign multm_ps2 = multm_reduce_add3b0_xor3b_wx2 ^ multm_reduce_sd2;
  assign multm_ps3 = multm_reduce_add3b0_xor3b_wx3 ^ multm_reduce_sd3;
  assign multm_ps4 = multm_reduce_add3b0_xor3b_wx4 ^ multm_reduce_sd4;
  assign multm_ps5 = multm_reduce_add3b0_xor3b_wx5 ^ multm_reduce_sd5;
  assign multm_ps6 = multm_reduce_add3b0_xor3b_wx6 ^ multm_reduce_sd6;
  assign multm_ps7 = multm_reduce_add3b0_xor3b_wx7 ^ multm_reduce_sd7;
  assign multm_ps8 = multm_reduce_add3b0_xor3b_wx8 ^ multm_reduce_sd8;
  assign multm_ps9 = multm_reduce_add3b0_xor3b_wx9 ^ multm_reduce_sd9;
  assign multm_ps10 = multm_reduce_add3b0_xor3b_wx10 ^ multm_reduce_sd10;
  assign multm_ps11 = multm_reduce_add3b1_xor3b_wx0 ^ multm_reduce_mc10;
  assign multm_ps12 = multm_reduce_add3b1_xor3b_wx1 ^ multm_reduce_mc11;
  assign multm_ps13 = multm_reduce_add3b1_xor3b_wx2 ^ multm_reduce_mc12;
  assign multm_ps14 = multm_reduce_add3b1_xor3b_wx3 ^ multm_reduce_mc13;
  assign multm_ps15 = multm_reduce_add3b1_xor3b_wx4 ^ multm_reduce_mc14;
  assign multm_ps16 = multm_reduce_add3b1_xor3b_wx5 ^ multm_reduce_mc15;
  assign multm_ps17 = multm_reduce_add3b1_xor3b_wx6 ^ multm_reduce_mc16;
  assign multm_ps18 = multm_reduce_add3b1_xor3b_wx7 ^ multm_reduce_mc17;
  assign multm_ps19 = multm_reduce_add3b1_xor3b_wx8 ^ multm_reduce_mc18;
  assign multm_ps20 = multm_reduce_add3b1_xor3b_wx9 ^ multm_reduce_mc19;
  assign multm_ps21 = multm_reduce_add3b1_xor3b_wx10 ^ multm_reduce_mc20;
  assign multm_ps22 = multm_reduce_add3b1_xor3b_wx11 ^ multm_reduce_mc21;
  assign multm_ps23 = multm_reduce_add3b1_xor3b_wx12 ^ multm_reduce_mc22;
  assign multm_ps24 = multm_reduce_add3b1_xor3b_wx13 ^ multm_reduce_mc23;
  assign multm_ps25 = multm_reduce_add3b1_xor3b_wx14 ^ multm_reduce_mc24;
  assign multm_ps26 = multm_reduce_add3b1_xor3b_wx15 ^ multm_reduce_mc25;
  assign multm_ps27 = multm_reduce_add3b1_xor3b_wx16 ^ multm_reduce_mc26;
  assign multm_ps28 = multm_reduce_add3b1_xor3b_wx17 ^ multm_reduce_mc27;
  assign multm_ps29 = multm_reduce_add3b1_xor3b_wx18 ^ multm_reduce_mc28;
  assign multm_ps30 = multm_reduce_add3b1_xor3b_wx19 ^ multm_reduce_mc29;
  assign multm_ps31 = multm_reduce_add3b1_xor3b_wx20 ^ multm_reduce_mc30;
  assign multm_ps32 = multm_reduce_add3b1_xor3b_wx21 ^ multm_reduce_mc31;
  assign multm_ps33 = multm_reduce_add3b1_xor3b_wx22 ^ multm_reduce_mc32;
  assign multm_ps34 = multm_reduce_add3b1_xor3b_wx23 ^ multm_reduce_mc33;
  assign multm_ps35 = multm_reduce_add3b1_xor3b_wx24 ^ multm_reduce_mc34;
  assign multm_ps36 = multm_reduce_add3b1_xor3b_wx25 ^ multm_reduce_mc35;
  assign multm_ps37 = multm_reduce_add3b1_xor3b_wx26 ^ multm_reduce_mc36;
  assign multm_ps38 = multm_reduce_add3b1_xor3b_wx27 ^ multm_reduce_mc37;
  assign multm_ps39 = multm_reduce_add3b1_xor3b_wx28 ^ multm_reduce_mc38;
  assign multm_ps40 = multm_reduce_add3b1_xor3b_wx29 ^ multm_reduce_mc39;
  assign multm_ps41 = multm_reduce_add3b1_xor3b_wx30 ^ multm_reduce_mc40;
  assign multm_ps42 = multm_reduce_add3b1_xor3b_wx31 ^ multm_reduce_mc41;
  assign multm_ps43 = multm_reduce_add3b1_xor3b_wx32 ^ multm_reduce_mc42;
  assign multm_ps44 = multm_reduce_add3b1_xor3b_wx33 ^ multm_reduce_mc43;
  assign multm_ps45 = multm_reduce_add3b1_xor3b_wx34 ^ multm_reduce_mc44;
  assign multm_ps46 = multm_reduce_add3b1_xor3b_wx35 ^ multm_reduce_mc45;
  assign multm_ps47 = multm_reduce_add3b1_xor3b_wx36 ^ multm_reduce_mc46;
  assign multm_ps48 = multm_reduce_add3b1_xor3b_wx37 ^ multm_reduce_mc47;
  assign multm_ps49 = multm_reduce_add3b1_xor3b_wx38 ^ multm_reduce_mc48;
  assign multm_ps50 = multm_reduce_add3b1_xor3b_wx39 ^ multm_reduce_mc49;
  assign multm_ps51 = multm_reduce_add3b1_xor3b_wx40 ^ multm_reduce_mc50;
  assign multm_ps52 = multm_reduce_add3b1_xor3b_wx41 ^ multm_reduce_mc51;
  assign multm_ps53 = multm_reduce_add3b1_xor3b_wx42 ^ multm_reduce_mc52;
  assign multm_ps54 = multm_reduce_add3b1_xor3b_wx43 ^ multm_reduce_mc53;
  assign multm_ps55 = multm_reduce_add3b1_xor3b_wx44 ^ multm_reduce_mc54;
  assign multm_ps56 = multm_reduce_add3b1_xor3b_wx45 ^ multm_reduce_mc55;
  assign multm_ps57 = multm_reduce_add3b1_xor3b_wx46 ^ multm_reduce_mc56;
  assign multm_ps58 = multm_reduce_add3b1_xor3b_wx47 ^ multm_reduce_mc57;
  assign multm_ps59 = multm_reduce_add3b1_xor3b_wx48 ^ multm_reduce_mc58;
  assign multm_ps60 = multm_reduce_add3b1_xor3b_wx49 ^ multm_reduce_mc59;
  assign multm_ps61 = multm_reduce_add3b1_xor3b_wx50 ^ multm_reduce_mc60;
  assign multm_ps62 = multm_reduce_add3b1_xor3b_wx51 ^ multm_reduce_mc61;
  assign multm_ps63 = multm_reduce_add3b1_xor3b_wx52 ^ multm_reduce_mc62;
  assign multm_ps64 = multm_reduce_add3b1_xor3b_wx53 ^ multm_reduce_mc63;
  assign multm_ps65 = multm_reduce_add3b1_xor3b_wx54 ^ multm_reduce_mc64;
  assign multm_ps66 = multm_reduce_add3b1_xor3b_wx55 ^ multm_reduce_mc65;
  assign multm_ps67 = multm_reduce_add3b1_xor3b_wx56 ^ multm_reduce_mc66;
  assign multm_ps68 = multm_reduce_add3b1_xor3b_wx57 ^ multm_reduce_mc67;
  assign multm_ps69 = multm_reduce_add3b1_xor3b_wx58 ^ multm_reduce_mc68;
  assign multm_ps70 = multm_reduce_add3b1_xor3b_wx59 ^ multm_reduce_mc69;
  assign multm_ps71 = multm_reduce_add3b1_xor3b_wx60 ^ multm_reduce_mc70;
  assign multm_ps72 = multm_reduce_add3b1_xor3b_wx61 ^ multm_reduce_mc71;
  assign multm_ps73 = multm_reduce_add3b1_xor3b_wx62 ^ multm_reduce_mc72;
  assign multm_ps74 = multm_reduce_add3b1_xor3b_wx63 ^ multm_reduce_mc73;
  assign multm_ps75 = multm_reduce_add3b1_xor3b_wx64 ^ multm_reduce_mc74;
  assign multm_ps76 = multm_reduce_add3b1_xor3b_wx65 ^ multm_reduce_mc75;
  assign multm_ps77 = multm_reduce_add3b1_xor3b_wx66 ^ multm_reduce_mc76;
  assign multm_ps78 = multm_reduce_add3b1_xor3b_wx67 ^ multm_reduce_mc77;
  assign multm_ps79 = multm_reduce_add3b1_xor3b_wx68 ^ multm_reduce_mc78;
  assign multm_ps80 = multm_reduce_add3b1_xor3b_wx69 ^ multm_reduce_mc79;
  assign multm_ps81 = multm_reduce_add3b1_xor3b_wx70 ^ multm_reduce_mc80;
  assign multm_ps82 = multm_reduce_add3b1_xor3b_wx71 ^ multm_reduce_mc81;
  assign multm_ps83 = multm_reduce_add3b1_xor3b_wx72 ^ multm_reduce_mc82;
  assign multm_ps84 = multm_reduce_add3b1_xor3b_wx73 ^ multm_reduce_mc83;
  assign multm_ps85 = multm_reduce_add3b1_xor3b_wx74 ^ multm_reduce_mc84;
  assign multm_ps86 = multm_reduce_add3b1_xor3b_wx75 ^ multm_reduce_mc85;
  assign multm_ps87 = multm_reduce_add3b1_xor3b_wx76 ^ multm_reduce_mc86;
  assign multm_ps88 = multm_reduce_add3b1_xor3b_wx77 ^ multm_reduce_mc87;
  assign multm_ps89 = multm_reduce_add3b1_xor3b_wx78 ^ multm_reduce_mc88;
  assign multm_ps90 = multm_reduce_add3b1_xor3b_wx79 ^ multm_reduce_mc89;
  assign multm_ps91 = multm_reduce_add3b1_xor3b_wx80 ^ multm_reduce_mc90;
  assign multm_ps92 = multm_reduce_add3b1_xor3b_wx81 ^ multm_reduce_mc91;
  assign multm_ps93 = multm_reduce_add3b1_xor3b_wx82 ^ multm_reduce_mc92;
  assign multm_ps94 = multm_reduce_add3b1_xor3b_wx83 ^ multm_reduce_mc93;
  assign multm_ps95 = multm_reduce_add3b1_xor3b_wx84 ^ multm_reduce_mc94;
  assign multm_ps96 = multm_reduce_add3b1_xor3b_wx85 ^ multm_reduce_mc95;
  assign multm_ps97 = multm_reduce_add3b1_xor3b_wx86 ^ multm_reduce_mc96;
  assign multm_ps98 = multm_reduce_add3b1_xor3b_wx87 ^ multm_reduce_mc97;
  assign multm_ps99 = multm_reduce_add3b1_xor3b_wx88 ^ multm_reduce_mc98;
  assign multm_ps100 = multm_reduce_add3b1_xor3b_wx89 ^ multm_reduce_mc99;
  assign multm_ps101 = multm_reduce_add3b1_xor3b_wx90 ^ multm_reduce_mc100;
  assign multm_ps102 = multm_reduce_add3b1_xor3b_wx91 ^ multm_reduce_mc101;
  assign multm_ps103 = multm_reduce_add3b1_xor3b_wx92 ^ multm_reduce_mc102;
  assign multm_ps104 = multm_reduce_add3b1_xor3b_wx93 ^ multm_reduce_mc103;
  assign multm_ps105 = multm_reduce_add3b1_xor3b_wx94 ^ multm_reduce_mc104;
  assign multm_ps106 = multm_reduce_add3b1_xor3b_wx95 ^ multm_reduce_mc105;
  assign multm_ps107 = multm_reduce_add3b1_xor3b_wx96 ^ multm_reduce_mc106;
  assign multm_ps108 = multm_reduce_add3b1_xor3b_wx97 ^ multm_reduce_mc107;
  assign multm_ps109 = multm_reduce_add3b1_xor3b_wx98 ^ multm_reduce_mc108;
  assign multm_ps110 = multm_reduce_add3b1_xor3b_wx99 ^ multm_reduce_mc109;
  assign multm_ps111 = multm_reduce_add3b1_xor3b_wx100 ^ multm_reduce_mc110;
  assign multm_ps112 = multm_reduce_add3b1_xor3b_wx101 ^ multm_reduce_mc111;
  assign multm_ps113 = multm_reduce_add3b1_xor3b_wx102 ^ multm_reduce_mc112;
  assign multm_ps114 = multm_reduce_add3b1_xor3b_wx103 ^ multm_reduce_mc113;
  assign multm_ps115 = multm_reduce_add3b1_xor3b_wx104 ^ multm_reduce_mc114;
  assign multm_ps116 = multm_reduce_add3b1_xor3b_wx105 ^ multm_reduce_mc115;
  assign multm_ps117 = multm_reduce_add3b1_xor3b_wx106 ^ multm_reduce_mc116;
  assign multm_ps118 = multm_reduce_add3b1_xor3b_wx107 ^ multm_reduce_mc117;
  assign multm_ps119 = multm_reduce_add3b1_xor3b_wx108 ^ multm_reduce_mc118;
  assign multm_ps120 = multm_reduce_add3b1_xor3b_wx109 ^ multm_reduce_mc119;
  assign multm_ps121 = multm_reduce_add3b1_xor3b_wx110 ^ multm_reduce_mc120;
  assign multm_ps122 = multm_reduce_add3b1_xor3b_wx111 ^ multm_reduce_mc121;
  assign multm_ps123 = multm_reduce_add3b1_xor3b_wx112 ^ multm_reduce_mc122;
  assign multm_ps124 = multm_reduce_add3b1_xor3b_wx113 ^ multm_reduce_mc123;
  assign multm_ps125 = multm_reduce_add3b1_xor3b_wx114 ^ multm_reduce_mc124;
  assign multm_ps126 = multm_reduce_add3b1_xor3b_wx115 ^ multm_reduce_mc125;
  assign multm_ps127 = multm_reduce_add3b1_xor3b_wx116 ^ multm_reduce_mc126;
  assign multm_ps128 = multm_reduce_add3b1_xor3b_wx117 ^ multm_reduce_mc127;
  assign multm_ps129 = multm_reduce_add3b1_xor3b_wx118 ^ multm_reduce_mc128;
  assign multm_ps130 = multm_reduce_add3b1_xor3b_wx119 ^ multm_reduce_mc129;
  assign multm_ps131 = multm_reduce_add3b1_xor3b_wx120 ^ multm_reduce_mc130;
  assign multm_ps132 = multm_reduce_add3b1_xor3b_wx121 ^ multm_reduce_mc131;
  assign multm_ps133 = multm_reduce_add3b1_xor3b_wx122 ^ multm_reduce_mc132;
  assign multm_ps134 = multm_reduce_add3b1_xor3b_wx123 ^ multm_reduce_mc133;
  assign multm_ps135 = multm_reduce_add3b1_xor3b_wx124 ^ multm_reduce_mc134;
  assign multm_ps136 = multm_reduce_add3b1_xor3b_wx125 ^ multm_reduce_mc135;
  assign multm_ps137 = multm_reduce_add3b1_xor3b_wx126 ^ multm_reduce_mc136;
  assign multm_ps138 = multm_reduce_add3b1_xor3b_wx127 ^ multm_reduce_mc137;
  assign multm_ps139 = multm_reduce_add3b1_xor3b_wx128 ^ multm_reduce_mc138;
  assign multm_ps140 = multm_reduce_add3b1_xor3b_wx129 ^ multm_reduce_mc139;
  assign multm_ps141 = multm_reduce_add3b1_xor3b_wx130 ^ multm_reduce_mc140;
  assign multm_ps142 = multm_reduce_add3b1_xor3b_wx131 ^ multm_reduce_mc141;
  assign multm_ps143 = multm_reduce_add3b1_xor3b_wx132 ^ multm_reduce_mc142;
  assign multm_ps144 = multm_reduce_add3b1_xor3b_wx133 ^ multm_reduce_mc143;
  assign multm_ps145 = multm_reduce_add3b1_xor3b_wx134 ^ multm_reduce_mc144;
  assign multm_ps146 = multm_reduce_add3b1_xor3b_wx135 ^ multm_reduce_mc145;
  assign multm_ps147 = multm_reduce_add3b1_xor3b_wx136 ^ multm_reduce_mc146;
  assign multm_ps148 = multm_reduce_add3b1_xor3b_wx137 ^ multm_reduce_mc147;
  assign multm_ps149 = multm_reduce_add3b1_xor3b_wx138 ^ multm_reduce_mc148;
  assign multm_ps150 = multm_reduce_add3b1_xor3b_wx139 ^ multm_reduce_mc149;
  assign multm_ps151 = multm_reduce_add3b1_xor3b_wx140 ^ multm_reduce_mc150;
  assign multm_ps152 = multm_reduce_add3b1_xor3b_wx141 ^ multm_reduce_mc151;
  assign multm_ps153 = multm_reduce_add3b1_xor3b_wx142 ^ multm_reduce_mc152;
  assign multm_ps154 = multm_reduce_add3b1_xor3b_wx143 ^ multm_reduce_mc153;
  assign multm_ps155 = multm_reduce_add3b1_xor3b_wx144 ^ multm_reduce_mc154;
  assign multm_ps156 = multm_reduce_add3b1_xor3b_wx145 ^ multm_reduce_mc155;
  assign multm_ps157 = multm_reduce_add3b1_xor3b_wx146 ^ multm_reduce_mc156;
  assign multm_ps158 = multm_reduce_add3b1_xor3b_wx147 ^ multm_reduce_mc157;
  assign multm_ps159 = multm_reduce_add3b1_xor3b_wx148 ^ multm_reduce_mc158;
  assign multm_ps160 = multm_reduce_add3b1_xor3b_wx149 ^ multm_reduce_mc159;
  assign multm_ps161 = multm_reduce_add3b1_xor3b_wx150 ^ multm_reduce_mc160;
  assign multm_ps162 = multm_reduce_add3b1_xor3b_wx151 ^ multm_reduce_mc161;
  assign multm_ps163 = multm_reduce_add3b1_xor3b_wx152 ^ multm_reduce_mc162;
  assign multm_ps164 = multm_reduce_add3b1_xor3b_wx153 ^ multm_reduce_mc163;
  assign multm_ps165 = multm_reduce_add3b1_xor3b_wx154 ^ multm_reduce_mc164;
  assign multm_ps166 = multm_reduce_add3b1_xor3b_wx155 ^ multm_reduce_mc165;
  assign multm_ps167 = multm_reduce_add3b1_xor3b_wx156 ^ multm_reduce_mc166;
  assign multm_ps168 = multm_reduce_add3b1_xor3b_wx157 ^ multm_reduce_mc167;
  assign multm_ps169 = multm_reduce_add3b1_xor3b_wx158 ^ multm_reduce_mc168;
  assign multm_ps170 = multm_reduce_add3b1_xor3b_wx159 ^ multm_reduce_mc169;
  assign multm_ps171 = multm_reduce_add3b1_xor3b_wx160 ^ multm_reduce_mc170;
  assign multm_ps172 = multm_reduce_add3b1_xor3b_wx161 ^ multm_reduce_mc171;
  assign multm_ps173 = multm_reduce_add3b1_xor3b_wx162 ^ multm_reduce_mc172;
  assign multm_ps174 = multm_reduce_add3b1_xor3b_wx163 ^ multm_reduce_mc173;
  assign multm_ps175 = multm_reduce_add3b1_xor3b_wx164 ^ multm_reduce_mc174;
  assign multm_ps176 = multm_reduce_add3b1_xor3b_wx165 ^ multm_reduce_mc175;
  assign multm_ps177 = multm_reduce_add3b1_xor3b_wx166 ^ multm_reduce_mc176;
  assign multm_ps178 = multm_reduce_add3b1_xor3b_wx167 ^ multm_reduce_mc177;
  assign multm_ps179 = multm_reduce_add3b1_xor3b_wx168 ^ multm_reduce_mc178;
  assign multm_ps180 = multm_reduce_add3b1_xor3b_wx169 ^ multm_reduce_mc179;
  assign multm_ps181 = multm_reduce_add3b1_xor3b_wx170 ^ multm_reduce_mc180;
  assign multm_ps182 = multm_reduce_add3b1_xor3b_wx171 ^ multm_reduce_mc181;
  assign multm_ps183 = multm_reduce_add3b1_xor3b_wx172 ^ multm_reduce_mc182;
  assign multm_ps184 = multm_reduce_add3_xor3_wx ^ multm_reduce_mc183;
  assign multm_qcr0 = multm_jpd ? multm_pc0 : multm_qcp0;
  assign multm_qcr1 = multm_jpd ? multm_pc1 : multm_qcp1;
  assign multm_qcr2 = multm_jpd ? multm_pc2 : multm_qcp2;
  assign multm_qcr3 = multm_jpd ? multm_pc3 : multm_qcp3;
  assign multm_qcr4 = multm_jpd ? multm_pc4 : multm_qcp4;
  assign multm_qcr5 = multm_jpd ? multm_pc5 : multm_qcp5;
  assign multm_qcr6 = multm_jpd ? multm_pc6 : multm_qcp6;
  assign multm_qcr7 = multm_jpd ? multm_pc7 : multm_qcp7;
  assign multm_qcr8 = multm_jpd ? multm_pc8 : multm_qcp8;
  assign multm_qcr9 = multm_jpd ? multm_pc9 : multm_qcp9;
  assign multm_qcr10 = xn0 & multm_qcp10;
  assign multm_qcr11 = multm_jpd ? multm_pc11 : multm_qcp11;
  assign multm_qcr12 = multm_jpd ? multm_pc12 : multm_qcp12;
  assign multm_qcr13 = multm_jpd ? multm_pc13 : multm_qcp13;
  assign multm_qcr14 = multm_jpd ? multm_pc14 : multm_qcp14;
  assign multm_qcr15 = multm_jpd ? multm_pc15 : multm_qcp15;
  assign multm_qcr16 = multm_jpd ? multm_pc16 : multm_qcp16;
  assign multm_qcr17 = multm_jpd ? multm_pc17 : multm_qcp17;
  assign multm_qcr18 = multm_jpd ? multm_pc18 : multm_qcp18;
  assign multm_qcr19 = multm_jpd ? multm_pc19 : multm_qcp19;
  assign multm_qcr20 = multm_jpd ? multm_pc20 : multm_qcp20;
  assign multm_qcr21 = multm_jpd ? multm_pc21 : multm_qcp21;
  assign multm_qcr22 = multm_jpd ? multm_pc22 : multm_qcp22;
  assign multm_qcr23 = multm_jpd ? multm_pc23 : multm_qcp23;
  assign multm_qcr24 = multm_jpd ? multm_pc24 : multm_qcp24;
  assign multm_qcr25 = multm_jpd ? multm_pc25 : multm_qcp25;
  assign multm_qcr26 = multm_jpd ? multm_pc26 : multm_qcp26;
  assign multm_qcr27 = multm_jpd ? multm_pc27 : multm_qcp27;
  assign multm_qcr28 = multm_jpd ? multm_pc28 : multm_qcp28;
  assign multm_qcr29 = multm_jpd ? multm_pc29 : multm_qcp29;
  assign multm_qcr30 = multm_jpd ? multm_pc30 : multm_qcp30;
  assign multm_qcr31 = multm_jpd ? multm_pc31 : multm_qcp31;
  assign multm_qcr32 = multm_jpd ? multm_pc32 : multm_qcp32;
  assign multm_qcr33 = multm_jpd ? multm_pc33 : multm_qcp33;
  assign multm_qcr34 = multm_jpd ? multm_pc34 : multm_qcp34;
  assign multm_qcr35 = multm_jpd ? multm_pc35 : multm_qcp35;
  assign multm_qcr36 = multm_jpd ? multm_pc36 : multm_qcp36;
  assign multm_qcr37 = multm_jpd ? multm_pc37 : multm_qcp37;
  assign multm_qcr38 = multm_jpd ? multm_pc38 : multm_qcp38;
  assign multm_qcr39 = multm_jpd ? multm_pc39 : multm_qcp39;
  assign multm_qcr40 = multm_jpd ? multm_pc40 : multm_qcp40;
  assign multm_qcr41 = multm_jpd ? multm_pc41 : multm_qcp41;
  assign multm_qcr42 = multm_jpd ? multm_pc42 : multm_qcp42;
  assign multm_qcr43 = multm_jpd ? multm_pc43 : multm_qcp43;
  assign multm_qcr44 = multm_jpd ? multm_pc44 : multm_qcp44;
  assign multm_qcr45 = multm_jpd ? multm_pc45 : multm_qcp45;
  assign multm_qcr46 = multm_jpd ? multm_pc46 : multm_qcp46;
  assign multm_qcr47 = multm_jpd ? multm_pc47 : multm_qcp47;
  assign multm_qcr48 = multm_jpd ? multm_pc48 : multm_qcp48;
  assign multm_qcr49 = multm_jpd ? multm_pc49 : multm_qcp49;
  assign multm_qcr50 = multm_jpd ? multm_pc50 : multm_qcp50;
  assign multm_qcr51 = multm_jpd ? multm_pc51 : multm_qcp51;
  assign multm_qcr52 = multm_jpd ? multm_pc52 : multm_qcp52;
  assign multm_qcr53 = multm_jpd ? multm_pc53 : multm_qcp53;
  assign multm_qcr54 = multm_jpd ? multm_pc54 : multm_qcp54;
  assign multm_qcr55 = multm_jpd ? multm_pc55 : multm_qcp55;
  assign multm_qcr56 = multm_jpd ? multm_pc56 : multm_qcp56;
  assign multm_qcr57 = multm_jpd ? multm_pc57 : multm_qcp57;
  assign multm_qcr58 = multm_jpd ? multm_pc58 : multm_qcp58;
  assign multm_qcr59 = multm_jpd ? multm_pc59 : multm_qcp59;
  assign multm_qcr60 = multm_jpd ? multm_pc60 : multm_qcp60;
  assign multm_qcr61 = multm_jpd ? multm_pc61 : multm_qcp61;
  assign multm_qcr62 = multm_jpd ? multm_pc62 : multm_qcp62;
  assign multm_qcr63 = multm_jpd ? multm_pc63 : multm_qcp63;
  assign multm_qcr64 = multm_jpd ? multm_pc64 : multm_qcp64;
  assign multm_qcr65 = multm_jpd ? multm_pc65 : multm_qcp65;
  assign multm_qcr66 = multm_jpd ? multm_pc66 : multm_qcp66;
  assign multm_qcr67 = multm_jpd ? multm_pc67 : multm_qcp67;
  assign multm_qcr68 = multm_jpd ? multm_pc68 : multm_qcp68;
  assign multm_qcr69 = multm_jpd ? multm_pc69 : multm_qcp69;
  assign multm_qcr70 = multm_jpd ? multm_pc70 : multm_qcp70;
  assign multm_qcr71 = multm_jpd ? multm_pc71 : multm_qcp71;
  assign multm_qcr72 = multm_jpd ? multm_pc72 : multm_qcp72;
  assign multm_qcr73 = multm_jpd ? multm_pc73 : multm_qcp73;
  assign multm_qcr74 = multm_jpd ? multm_pc74 : multm_qcp74;
  assign multm_qcr75 = multm_jpd ? multm_pc75 : multm_qcp75;
  assign multm_qcr76 = multm_jpd ? multm_pc76 : multm_qcp76;
  assign multm_qcr77 = multm_jpd ? multm_pc77 : multm_qcp77;
  assign multm_qcr78 = multm_jpd ? multm_pc78 : multm_qcp78;
  assign multm_qcr79 = multm_jpd ? multm_pc79 : multm_qcp79;
  assign multm_qcr80 = multm_jpd ? multm_pc80 : multm_qcp80;
  assign multm_qcr81 = multm_jpd ? multm_pc81 : multm_qcp81;
  assign multm_qcr82 = multm_jpd ? multm_pc82 : multm_qcp82;
  assign multm_qcr83 = multm_jpd ? multm_pc83 : multm_qcp83;
  assign multm_qcr84 = multm_jpd ? multm_pc84 : multm_qcp84;
  assign multm_qcr85 = multm_jpd ? multm_pc85 : multm_qcp85;
  assign multm_qcr86 = multm_jpd ? multm_pc86 : multm_qcp86;
  assign multm_qcr87 = multm_jpd ? multm_pc87 : multm_qcp87;
  assign multm_qcr88 = multm_jpd ? multm_pc88 : multm_qcp88;
  assign multm_qcr89 = multm_jpd ? multm_pc89 : multm_qcp89;
  assign multm_qcr90 = multm_jpd ? multm_pc90 : multm_qcp90;
  assign multm_qcr91 = multm_jpd ? multm_pc91 : multm_qcp91;
  assign multm_qcr92 = multm_jpd ? multm_pc92 : multm_qcp92;
  assign multm_qcr93 = multm_jpd ? multm_pc93 : multm_qcp93;
  assign multm_qcr94 = multm_jpd ? multm_pc94 : multm_qcp94;
  assign multm_qcr95 = multm_jpd ? multm_pc95 : multm_qcp95;
  assign multm_qcr96 = multm_jpd ? multm_pc96 : multm_qcp96;
  assign multm_qcr97 = multm_jpd ? multm_pc97 : multm_qcp97;
  assign multm_qcr98 = multm_jpd ? multm_pc98 : multm_qcp98;
  assign multm_qcr99 = multm_jpd ? multm_pc99 : multm_qcp99;
  assign multm_qcr100 = multm_jpd ? multm_pc100 : multm_qcp100;
  assign multm_qcr101 = multm_jpd ? multm_pc101 : multm_qcp101;
  assign multm_qcr102 = multm_jpd ? multm_pc102 : multm_qcp102;
  assign multm_qcr103 = multm_jpd ? multm_pc103 : multm_qcp103;
  assign multm_qcr104 = multm_jpd ? multm_pc104 : multm_qcp104;
  assign multm_qcr105 = multm_jpd ? multm_pc105 : multm_qcp105;
  assign multm_qcr106 = multm_jpd ? multm_pc106 : multm_qcp106;
  assign multm_qcr107 = multm_jpd ? multm_pc107 : multm_qcp107;
  assign multm_qcr108 = multm_jpd ? multm_pc108 : multm_qcp108;
  assign multm_qcr109 = multm_jpd ? multm_pc109 : multm_qcp109;
  assign multm_qcr110 = multm_jpd ? multm_pc110 : multm_qcp110;
  assign multm_qcr111 = multm_jpd ? multm_pc111 : multm_qcp111;
  assign multm_qcr112 = multm_jpd ? multm_pc112 : multm_qcp112;
  assign multm_qcr113 = multm_jpd ? multm_pc113 : multm_qcp113;
  assign multm_qcr114 = multm_jpd ? multm_pc114 : multm_qcp114;
  assign multm_qcr115 = multm_jpd ? multm_pc115 : multm_qcp115;
  assign multm_qcr116 = multm_jpd ? multm_pc116 : multm_qcp116;
  assign multm_qcr117 = multm_jpd ? multm_pc117 : multm_qcp117;
  assign multm_qcr118 = multm_jpd ? multm_pc118 : multm_qcp118;
  assign multm_qcr119 = multm_jpd ? multm_pc119 : multm_qcp119;
  assign multm_qcr120 = multm_jpd ? multm_pc120 : multm_qcp120;
  assign multm_qcr121 = multm_jpd ? multm_pc121 : multm_qcp121;
  assign multm_qcr122 = multm_jpd ? multm_pc122 : multm_qcp122;
  assign multm_qcr123 = multm_jpd ? multm_pc123 : multm_qcp123;
  assign multm_qcr124 = multm_jpd ? multm_pc124 : multm_qcp124;
  assign multm_qcr125 = multm_jpd ? multm_pc125 : multm_qcp125;
  assign multm_qcr126 = multm_jpd ? multm_pc126 : multm_qcp126;
  assign multm_qcr127 = multm_jpd ? multm_pc127 : multm_qcp127;
  assign multm_qcr128 = multm_jpd ? multm_pc128 : multm_qcp128;
  assign multm_qcr129 = multm_jpd ? multm_pc129 : multm_qcp129;
  assign multm_qcr130 = multm_jpd ? multm_pc130 : multm_qcp130;
  assign multm_qcr131 = multm_jpd ? multm_pc131 : multm_qcp131;
  assign multm_qcr132 = multm_jpd ? multm_pc132 : multm_qcp132;
  assign multm_qcr133 = multm_jpd ? multm_pc133 : multm_qcp133;
  assign multm_qcr134 = multm_jpd ? multm_pc134 : multm_qcp134;
  assign multm_qcr135 = multm_jpd ? multm_pc135 : multm_qcp135;
  assign multm_qcr136 = multm_jpd ? multm_pc136 : multm_qcp136;
  assign multm_qcr137 = multm_jpd ? multm_pc137 : multm_qcp137;
  assign multm_qcr138 = multm_jpd ? multm_pc138 : multm_qcp138;
  assign multm_qcr139 = multm_jpd ? multm_pc139 : multm_qcp139;
  assign multm_qcr140 = multm_jpd ? multm_pc140 : multm_qcp140;
  assign multm_qcr141 = multm_jpd ? multm_pc141 : multm_qcp141;
  assign multm_qcr142 = multm_jpd ? multm_pc142 : multm_qcp142;
  assign multm_qcr143 = multm_jpd ? multm_pc143 : multm_qcp143;
  assign multm_qcr144 = multm_jpd ? multm_pc144 : multm_qcp144;
  assign multm_qcr145 = multm_jpd ? multm_pc145 : multm_qcp145;
  assign multm_qcr146 = multm_jpd ? multm_pc146 : multm_qcp146;
  assign multm_qcr147 = multm_jpd ? multm_pc147 : multm_qcp147;
  assign multm_qcr148 = multm_jpd ? multm_pc148 : multm_qcp148;
  assign multm_qcr149 = multm_jpd ? multm_pc149 : multm_qcp149;
  assign multm_qcr150 = multm_jpd ? multm_pc150 : multm_qcp150;
  assign multm_qcr151 = multm_jpd ? multm_pc151 : multm_qcp151;
  assign multm_qcr152 = multm_jpd ? multm_pc152 : multm_qcp152;
  assign multm_qcr153 = multm_jpd ? multm_pc153 : multm_qcp153;
  assign multm_qcr154 = multm_jpd ? multm_pc154 : multm_qcp154;
  assign multm_qcr155 = multm_jpd ? multm_pc155 : multm_qcp155;
  assign multm_qcr156 = multm_jpd ? multm_pc156 : multm_qcp156;
  assign multm_qcr157 = multm_jpd ? multm_pc157 : multm_qcp157;
  assign multm_qcr158 = multm_jpd ? multm_pc158 : multm_qcp158;
  assign multm_qcr159 = multm_jpd ? multm_pc159 : multm_qcp159;
  assign multm_qcr160 = multm_jpd ? multm_pc160 : multm_qcp160;
  assign multm_qcr161 = multm_jpd ? multm_pc161 : multm_qcp161;
  assign multm_qcr162 = multm_jpd ? multm_pc162 : multm_qcp162;
  assign multm_qcr163 = multm_jpd ? multm_pc163 : multm_qcp163;
  assign multm_qcr164 = multm_jpd ? multm_pc164 : multm_qcp164;
  assign multm_qcr165 = multm_jpd ? multm_pc165 : multm_qcp165;
  assign multm_qcr166 = multm_jpd ? multm_pc166 : multm_qcp166;
  assign multm_qcr167 = multm_jpd ? multm_pc167 : multm_qcp167;
  assign multm_qcr168 = multm_jpd ? multm_pc168 : multm_qcp168;
  assign multm_qcr169 = multm_jpd ? multm_pc169 : multm_qcp169;
  assign multm_qcr170 = multm_jpd ? multm_pc170 : multm_qcp170;
  assign multm_qcr171 = multm_jpd ? multm_pc171 : multm_qcp171;
  assign multm_qcr172 = multm_jpd ? multm_pc172 : multm_qcp172;
  assign multm_qcr173 = multm_jpd ? multm_pc173 : multm_qcp173;
  assign multm_qcr174 = multm_jpd ? multm_pc174 : multm_qcp174;
  assign multm_qcr175 = multm_jpd ? multm_pc175 : multm_qcp175;
  assign multm_qcr176 = multm_jpd ? multm_pc176 : multm_qcp176;
  assign multm_qcr177 = multm_jpd ? multm_pc177 : multm_qcp177;
  assign multm_qcr178 = multm_jpd ? multm_pc178 : multm_qcp178;
  assign multm_qcr179 = multm_jpd ? multm_pc179 : multm_qcp179;
  assign multm_qcr180 = multm_jpd ? multm_pc180 : multm_qcp180;
  assign multm_qcr181 = multm_jpd ? multm_pc181 : multm_qcp181;
  assign multm_qcr182 = multm_jpd ? multm_pc182 : multm_qcp182;
  assign multm_qcr183 = multm_jpd ? multm_pc183 : multm_qcp183;
  assign multm_qcr184 = multm_jpd ? multm_pc184 : multm_qcp184;
  assign multm_qsr0 = multm_jpd ? multm_ps0 : multm_qsp0;
  assign multm_qsr1 = multm_jpd ? multm_ps1 : multm_qsp1;
  assign multm_qsr2 = multm_jpd ? multm_ps2 : multm_qsp2;
  assign multm_qsr3 = multm_jpd ? multm_ps3 : multm_qsp3;
  assign multm_qsr4 = multm_jpd ? multm_ps4 : multm_qsp4;
  assign multm_qsr5 = multm_jpd ? multm_ps5 : multm_qsp5;
  assign multm_qsr6 = multm_jpd ? multm_ps6 : multm_qsp6;
  assign multm_qsr7 = multm_jpd ? multm_ps7 : multm_qsp7;
  assign multm_qsr8 = multm_jpd ? multm_ps8 : multm_qsp8;
  assign multm_qsr9 = multm_jpd ? multm_ps9 : multm_qsp9;
  assign multm_qsr10 = multm_jpd ? multm_ps10 : multm_qsp10;
  assign multm_qsr11 = multm_jpd ? multm_ps11 : multm_qsp11;
  assign multm_qsr12 = multm_jpd ? multm_ps12 : multm_qsp12;
  assign multm_qsr13 = multm_jpd ? multm_ps13 : multm_qsp13;
  assign multm_qsr14 = multm_jpd ? multm_ps14 : multm_qsp14;
  assign multm_qsr15 = multm_jpd ? multm_ps15 : multm_qsp15;
  assign multm_qsr16 = multm_jpd ? multm_ps16 : multm_qsp16;
  assign multm_qsr17 = multm_jpd ? multm_ps17 : multm_qsp17;
  assign multm_qsr18 = multm_jpd ? multm_ps18 : multm_qsp18;
  assign multm_qsr19 = multm_jpd ? multm_ps19 : multm_qsp19;
  assign multm_qsr20 = multm_jpd ? multm_ps20 : multm_qsp20;
  assign multm_qsr21 = multm_jpd ? multm_ps21 : multm_qsp21;
  assign multm_qsr22 = multm_jpd ? multm_ps22 : multm_qsp22;
  assign multm_qsr23 = multm_jpd ? multm_ps23 : multm_qsp23;
  assign multm_qsr24 = multm_jpd ? multm_ps24 : multm_qsp24;
  assign multm_qsr25 = multm_jpd ? multm_ps25 : multm_qsp25;
  assign multm_qsr26 = multm_jpd ? multm_ps26 : multm_qsp26;
  assign multm_qsr27 = multm_jpd ? multm_ps27 : multm_qsp27;
  assign multm_qsr28 = multm_jpd ? multm_ps28 : multm_qsp28;
  assign multm_qsr29 = multm_jpd ? multm_ps29 : multm_qsp29;
  assign multm_qsr30 = multm_jpd ? multm_ps30 : multm_qsp30;
  assign multm_qsr31 = multm_jpd ? multm_ps31 : multm_qsp31;
  assign multm_qsr32 = multm_jpd ? multm_ps32 : multm_qsp32;
  assign multm_qsr33 = multm_jpd ? multm_ps33 : multm_qsp33;
  assign multm_qsr34 = multm_jpd ? multm_ps34 : multm_qsp34;
  assign multm_qsr35 = multm_jpd ? multm_ps35 : multm_qsp35;
  assign multm_qsr36 = multm_jpd ? multm_ps36 : multm_qsp36;
  assign multm_qsr37 = multm_jpd ? multm_ps37 : multm_qsp37;
  assign multm_qsr38 = multm_jpd ? multm_ps38 : multm_qsp38;
  assign multm_qsr39 = multm_jpd ? multm_ps39 : multm_qsp39;
  assign multm_qsr40 = multm_jpd ? multm_ps40 : multm_qsp40;
  assign multm_qsr41 = multm_jpd ? multm_ps41 : multm_qsp41;
  assign multm_qsr42 = multm_jpd ? multm_ps42 : multm_qsp42;
  assign multm_qsr43 = multm_jpd ? multm_ps43 : multm_qsp43;
  assign multm_qsr44 = multm_jpd ? multm_ps44 : multm_qsp44;
  assign multm_qsr45 = multm_jpd ? multm_ps45 : multm_qsp45;
  assign multm_qsr46 = multm_jpd ? multm_ps46 : multm_qsp46;
  assign multm_qsr47 = multm_jpd ? multm_ps47 : multm_qsp47;
  assign multm_qsr48 = multm_jpd ? multm_ps48 : multm_qsp48;
  assign multm_qsr49 = multm_jpd ? multm_ps49 : multm_qsp49;
  assign multm_qsr50 = multm_jpd ? multm_ps50 : multm_qsp50;
  assign multm_qsr51 = multm_jpd ? multm_ps51 : multm_qsp51;
  assign multm_qsr52 = multm_jpd ? multm_ps52 : multm_qsp52;
  assign multm_qsr53 = multm_jpd ? multm_ps53 : multm_qsp53;
  assign multm_qsr54 = multm_jpd ? multm_ps54 : multm_qsp54;
  assign multm_qsr55 = multm_jpd ? multm_ps55 : multm_qsp55;
  assign multm_qsr56 = multm_jpd ? multm_ps56 : multm_qsp56;
  assign multm_qsr57 = multm_jpd ? multm_ps57 : multm_qsp57;
  assign multm_qsr58 = multm_jpd ? multm_ps58 : multm_qsp58;
  assign multm_qsr59 = multm_jpd ? multm_ps59 : multm_qsp59;
  assign multm_qsr60 = multm_jpd ? multm_ps60 : multm_qsp60;
  assign multm_qsr61 = multm_jpd ? multm_ps61 : multm_qsp61;
  assign multm_qsr62 = multm_jpd ? multm_ps62 : multm_qsp62;
  assign multm_qsr63 = multm_jpd ? multm_ps63 : multm_qsp63;
  assign multm_qsr64 = multm_jpd ? multm_ps64 : multm_qsp64;
  assign multm_qsr65 = multm_jpd ? multm_ps65 : multm_qsp65;
  assign multm_qsr66 = multm_jpd ? multm_ps66 : multm_qsp66;
  assign multm_qsr67 = multm_jpd ? multm_ps67 : multm_qsp67;
  assign multm_qsr68 = multm_jpd ? multm_ps68 : multm_qsp68;
  assign multm_qsr69 = multm_jpd ? multm_ps69 : multm_qsp69;
  assign multm_qsr70 = multm_jpd ? multm_ps70 : multm_qsp70;
  assign multm_qsr71 = multm_jpd ? multm_ps71 : multm_qsp71;
  assign multm_qsr72 = multm_jpd ? multm_ps72 : multm_qsp72;
  assign multm_qsr73 = multm_jpd ? multm_ps73 : multm_qsp73;
  assign multm_qsr74 = multm_jpd ? multm_ps74 : multm_qsp74;
  assign multm_qsr75 = multm_jpd ? multm_ps75 : multm_qsp75;
  assign multm_qsr76 = multm_jpd ? multm_ps76 : multm_qsp76;
  assign multm_qsr77 = multm_jpd ? multm_ps77 : multm_qsp77;
  assign multm_qsr78 = multm_jpd ? multm_ps78 : multm_qsp78;
  assign multm_qsr79 = multm_jpd ? multm_ps79 : multm_qsp79;
  assign multm_qsr80 = multm_jpd ? multm_ps80 : multm_qsp80;
  assign multm_qsr81 = multm_jpd ? multm_ps81 : multm_qsp81;
  assign multm_qsr82 = multm_jpd ? multm_ps82 : multm_qsp82;
  assign multm_qsr83 = multm_jpd ? multm_ps83 : multm_qsp83;
  assign multm_qsr84 = multm_jpd ? multm_ps84 : multm_qsp84;
  assign multm_qsr85 = multm_jpd ? multm_ps85 : multm_qsp85;
  assign multm_qsr86 = multm_jpd ? multm_ps86 : multm_qsp86;
  assign multm_qsr87 = multm_jpd ? multm_ps87 : multm_qsp87;
  assign multm_qsr88 = multm_jpd ? multm_ps88 : multm_qsp88;
  assign multm_qsr89 = multm_jpd ? multm_ps89 : multm_qsp89;
  assign multm_qsr90 = multm_jpd ? multm_ps90 : multm_qsp90;
  assign multm_qsr91 = multm_jpd ? multm_ps91 : multm_qsp91;
  assign multm_qsr92 = multm_jpd ? multm_ps92 : multm_qsp92;
  assign multm_qsr93 = multm_jpd ? multm_ps93 : multm_qsp93;
  assign multm_qsr94 = multm_jpd ? multm_ps94 : multm_qsp94;
  assign multm_qsr95 = multm_jpd ? multm_ps95 : multm_qsp95;
  assign multm_qsr96 = multm_jpd ? multm_ps96 : multm_qsp96;
  assign multm_qsr97 = multm_jpd ? multm_ps97 : multm_qsp97;
  assign multm_qsr98 = multm_jpd ? multm_ps98 : multm_qsp98;
  assign multm_qsr99 = multm_jpd ? multm_ps99 : multm_qsp99;
  assign multm_qsr100 = multm_jpd ? multm_ps100 : multm_qsp100;
  assign multm_qsr101 = multm_jpd ? multm_ps101 : multm_qsp101;
  assign multm_qsr102 = multm_jpd ? multm_ps102 : multm_qsp102;
  assign multm_qsr103 = multm_jpd ? multm_ps103 : multm_qsp103;
  assign multm_qsr104 = multm_jpd ? multm_ps104 : multm_qsp104;
  assign multm_qsr105 = multm_jpd ? multm_ps105 : multm_qsp105;
  assign multm_qsr106 = multm_jpd ? multm_ps106 : multm_qsp106;
  assign multm_qsr107 = multm_jpd ? multm_ps107 : multm_qsp107;
  assign multm_qsr108 = multm_jpd ? multm_ps108 : multm_qsp108;
  assign multm_qsr109 = multm_jpd ? multm_ps109 : multm_qsp109;
  assign multm_qsr110 = multm_jpd ? multm_ps110 : multm_qsp110;
  assign multm_qsr111 = multm_jpd ? multm_ps111 : multm_qsp111;
  assign multm_qsr112 = multm_jpd ? multm_ps112 : multm_qsp112;
  assign multm_qsr113 = multm_jpd ? multm_ps113 : multm_qsp113;
  assign multm_qsr114 = multm_jpd ? multm_ps114 : multm_qsp114;
  assign multm_qsr115 = multm_jpd ? multm_ps115 : multm_qsp115;
  assign multm_qsr116 = multm_jpd ? multm_ps116 : multm_qsp116;
  assign multm_qsr117 = multm_jpd ? multm_ps117 : multm_qsp117;
  assign multm_qsr118 = multm_jpd ? multm_ps118 : multm_qsp118;
  assign multm_qsr119 = multm_jpd ? multm_ps119 : multm_qsp119;
  assign multm_qsr120 = multm_jpd ? multm_ps120 : multm_qsp120;
  assign multm_qsr121 = multm_jpd ? multm_ps121 : multm_qsp121;
  assign multm_qsr122 = multm_jpd ? multm_ps122 : multm_qsp122;
  assign multm_qsr123 = multm_jpd ? multm_ps123 : multm_qsp123;
  assign multm_qsr124 = multm_jpd ? multm_ps124 : multm_qsp124;
  assign multm_qsr125 = multm_jpd ? multm_ps125 : multm_qsp125;
  assign multm_qsr126 = multm_jpd ? multm_ps126 : multm_qsp126;
  assign multm_qsr127 = multm_jpd ? multm_ps127 : multm_qsp127;
  assign multm_qsr128 = multm_jpd ? multm_ps128 : multm_qsp128;
  assign multm_qsr129 = multm_jpd ? multm_ps129 : multm_qsp129;
  assign multm_qsr130 = multm_jpd ? multm_ps130 : multm_qsp130;
  assign multm_qsr131 = multm_jpd ? multm_ps131 : multm_qsp131;
  assign multm_qsr132 = multm_jpd ? multm_ps132 : multm_qsp132;
  assign multm_qsr133 = multm_jpd ? multm_ps133 : multm_qsp133;
  assign multm_qsr134 = multm_jpd ? multm_ps134 : multm_qsp134;
  assign multm_qsr135 = multm_jpd ? multm_ps135 : multm_qsp135;
  assign multm_qsr136 = multm_jpd ? multm_ps136 : multm_qsp136;
  assign multm_qsr137 = multm_jpd ? multm_ps137 : multm_qsp137;
  assign multm_qsr138 = multm_jpd ? multm_ps138 : multm_qsp138;
  assign multm_qsr139 = multm_jpd ? multm_ps139 : multm_qsp139;
  assign multm_qsr140 = multm_jpd ? multm_ps140 : multm_qsp140;
  assign multm_qsr141 = multm_jpd ? multm_ps141 : multm_qsp141;
  assign multm_qsr142 = multm_jpd ? multm_ps142 : multm_qsp142;
  assign multm_qsr143 = multm_jpd ? multm_ps143 : multm_qsp143;
  assign multm_qsr144 = multm_jpd ? multm_ps144 : multm_qsp144;
  assign multm_qsr145 = multm_jpd ? multm_ps145 : multm_qsp145;
  assign multm_qsr146 = multm_jpd ? multm_ps146 : multm_qsp146;
  assign multm_qsr147 = multm_jpd ? multm_ps147 : multm_qsp147;
  assign multm_qsr148 = multm_jpd ? multm_ps148 : multm_qsp148;
  assign multm_qsr149 = multm_jpd ? multm_ps149 : multm_qsp149;
  assign multm_qsr150 = multm_jpd ? multm_ps150 : multm_qsp150;
  assign multm_qsr151 = multm_jpd ? multm_ps151 : multm_qsp151;
  assign multm_qsr152 = multm_jpd ? multm_ps152 : multm_qsp152;
  assign multm_qsr153 = multm_jpd ? multm_ps153 : multm_qsp153;
  assign multm_qsr154 = multm_jpd ? multm_ps154 : multm_qsp154;
  assign multm_qsr155 = multm_jpd ? multm_ps155 : multm_qsp155;
  assign multm_qsr156 = multm_jpd ? multm_ps156 : multm_qsp156;
  assign multm_qsr157 = multm_jpd ? multm_ps157 : multm_qsp157;
  assign multm_qsr158 = multm_jpd ? multm_ps158 : multm_qsp158;
  assign multm_qsr159 = multm_jpd ? multm_ps159 : multm_qsp159;
  assign multm_qsr160 = multm_jpd ? multm_ps160 : multm_qsp160;
  assign multm_qsr161 = multm_jpd ? multm_ps161 : multm_qsp161;
  assign multm_qsr162 = multm_jpd ? multm_ps162 : multm_qsp162;
  assign multm_qsr163 = multm_jpd ? multm_ps163 : multm_qsp163;
  assign multm_qsr164 = multm_jpd ? multm_ps164 : multm_qsp164;
  assign multm_qsr165 = multm_jpd ? multm_ps165 : multm_qsp165;
  assign multm_qsr166 = multm_jpd ? multm_ps166 : multm_qsp166;
  assign multm_qsr167 = multm_jpd ? multm_ps167 : multm_qsp167;
  assign multm_qsr168 = multm_jpd ? multm_ps168 : multm_qsp168;
  assign multm_qsr169 = multm_jpd ? multm_ps169 : multm_qsp169;
  assign multm_qsr170 = multm_jpd ? multm_ps170 : multm_qsp170;
  assign multm_qsr171 = multm_jpd ? multm_ps171 : multm_qsp171;
  assign multm_qsr172 = multm_jpd ? multm_ps172 : multm_qsp172;
  assign multm_qsr173 = multm_jpd ? multm_ps173 : multm_qsp173;
  assign multm_qsr174 = multm_jpd ? multm_ps174 : multm_qsp174;
  assign multm_qsr175 = multm_jpd ? multm_ps175 : multm_qsp175;
  assign multm_qsr176 = multm_jpd ? multm_ps176 : multm_qsp176;
  assign multm_qsr177 = multm_jpd ? multm_ps177 : multm_qsp177;
  assign multm_qsr178 = multm_jpd ? multm_ps178 : multm_qsp178;
  assign multm_qsr179 = multm_jpd ? multm_ps179 : multm_qsp179;
  assign multm_qsr180 = multm_jpd ? multm_ps180 : multm_qsp180;
  assign multm_qsr181 = multm_jpd ? multm_ps181 : multm_qsp181;
  assign multm_qsr182 = multm_jpd ? multm_ps182 : multm_qsp182;
  assign multm_qsr183 = multm_jpd ? multm_ps183 : multm_qsp183;
  assign multm_qsr184 = multm_jpd ? multm_ps184 : multm_qsp184;
  assign multm_reduce_add3_maj3_or3_wx = multm_reduce_add3_maj3_wx | multm_reduce_add3_maj3_wy;
  assign multm_reduce_add3_maj3_wx = multm_reduce_sb173 & multm_reduce_sa184;
  assign multm_reduce_add3_maj3_wy = multm_reduce_sb173 & multm_reduce_mc183;
  assign multm_reduce_add3_maj3_xy = multm_reduce_sa184 & multm_reduce_mc183;
  assign multm_reduce_add3_xor3_wx = multm_reduce_sb173 ^ multm_reduce_sa184;
  assign multm_reduce_add3b0_maj3b_or3b_wx0 = multm_reduce_add3b0_maj3b_wx0 | multm_reduce_add3b0_maj3b_wy0;
  assign multm_reduce_add3b0_maj3b_or3b_wx1 = multm_reduce_add3b0_maj3b_wx1 | multm_reduce_add3b0_maj3b_wy1;
  assign multm_reduce_add3b0_maj3b_or3b_wx2 = multm_reduce_add3b0_maj3b_wx2 | multm_reduce_add3b0_maj3b_wy2;
  assign multm_reduce_add3b0_maj3b_or3b_wx3 = multm_reduce_add3b0_maj3b_wx3 | multm_reduce_add3b0_maj3b_wy3;
  assign multm_reduce_add3b0_maj3b_or3b_wx4 = multm_reduce_add3b0_maj3b_wx4 | multm_reduce_add3b0_maj3b_wy4;
  assign multm_reduce_add3b0_maj3b_or3b_wx5 = multm_reduce_add3b0_maj3b_wx5 | multm_reduce_add3b0_maj3b_wy5;
  assign multm_reduce_add3b0_maj3b_or3b_wx6 = multm_reduce_add3b0_maj3b_wx6 | multm_reduce_add3b0_maj3b_wy6;
  assign multm_reduce_add3b0_maj3b_or3b_wx7 = multm_reduce_add3b0_maj3b_wx7 | multm_reduce_add3b0_maj3b_wy7;
  assign multm_reduce_add3b0_maj3b_or3b_wx8 = multm_reduce_add3b0_maj3b_wx8 | multm_reduce_add3b0_maj3b_wy8;
  assign multm_reduce_add3b0_maj3b_or3b_wx9 = multm_reduce_add3b0_maj3b_wx9 | multm_reduce_add3b0_maj3b_wy9;
  assign multm_reduce_add3b0_maj3b_or3b_wx10 = multm_reduce_add3b0_maj3b_wx10 | multm_reduce_add3b0_maj3b_wy10;
  assign multm_reduce_add3b0_maj3b_or3b_wx11 = multm_reduce_add3b0_maj3b_wx11 | multm_reduce_add3b0_maj3b_wy11;
  assign multm_reduce_add3b0_maj3b_or3b_wx12 = multm_reduce_add3b0_maj3b_wx12 | multm_reduce_add3b0_maj3b_wy12;
  assign multm_reduce_add3b0_maj3b_or3b_wx13 = multm_reduce_add3b0_maj3b_wx13 | multm_reduce_add3b0_maj3b_wy13;
  assign multm_reduce_add3b0_maj3b_or3b_wx14 = multm_reduce_add3b0_maj3b_wx14 | multm_reduce_add3b0_maj3b_wy14;
  assign multm_reduce_add3b0_maj3b_or3b_wx15 = multm_reduce_add3b0_maj3b_wx15 | multm_reduce_add3b0_maj3b_wy15;
  assign multm_reduce_add3b0_maj3b_or3b_wx16 = multm_reduce_add3b0_maj3b_wx16 | multm_reduce_add3b0_maj3b_wy16;
  assign multm_reduce_add3b0_maj3b_or3b_wx17 = multm_reduce_add3b0_maj3b_wx17 | multm_reduce_add3b0_maj3b_wy17;
  assign multm_reduce_add3b0_maj3b_or3b_wx18 = multm_reduce_add3b0_maj3b_wx18 | multm_reduce_add3b0_maj3b_wy18;
  assign multm_reduce_add3b0_maj3b_or3b_wx19 = multm_reduce_add3b0_maj3b_wx19 | multm_reduce_add3b0_maj3b_wy19;
  assign multm_reduce_add3b0_maj3b_or3b_wx20 = multm_reduce_add3b0_maj3b_wx20 | multm_reduce_add3b0_maj3b_wy20;
  assign multm_reduce_add3b0_maj3b_or3b_wx21 = multm_reduce_add3b0_maj3b_wx21 | multm_reduce_add3b0_maj3b_wy21;
  assign multm_reduce_add3b0_maj3b_or3b_wx22 = multm_reduce_add3b0_maj3b_wx22 | multm_reduce_add3b0_maj3b_wy22;
  assign multm_reduce_add3b0_maj3b_or3b_wx23 = multm_reduce_add3b0_maj3b_wx23 | multm_reduce_add3b0_maj3b_wy23;
  assign multm_reduce_add3b0_maj3b_or3b_wx24 = multm_reduce_add3b0_maj3b_wx24 | multm_reduce_add3b0_maj3b_wy24;
  assign multm_reduce_add3b0_maj3b_or3b_wx25 = multm_reduce_add3b0_maj3b_wx25 | multm_reduce_add3b0_maj3b_wy25;
  assign multm_reduce_add3b0_maj3b_or3b_wx26 = multm_reduce_add3b0_maj3b_wx26 | multm_reduce_add3b0_maj3b_wy26;
  assign multm_reduce_add3b0_maj3b_or3b_wx27 = multm_reduce_add3b0_maj3b_wx27 | multm_reduce_add3b0_maj3b_wy27;
  assign multm_reduce_add3b0_maj3b_or3b_wx28 = multm_reduce_add3b0_maj3b_wx28 | multm_reduce_add3b0_maj3b_wy28;
  assign multm_reduce_add3b0_maj3b_or3b_wx29 = multm_reduce_add3b0_maj3b_wx29 | multm_reduce_add3b0_maj3b_wy29;
  assign multm_reduce_add3b0_maj3b_or3b_wx30 = multm_reduce_add3b0_maj3b_wx30 | multm_reduce_add3b0_maj3b_wy30;
  assign multm_reduce_add3b0_maj3b_or3b_wx31 = multm_reduce_add3b0_maj3b_wx31 | multm_reduce_add3b0_maj3b_wy31;
  assign multm_reduce_add3b0_maj3b_or3b_wx32 = multm_reduce_add3b0_maj3b_wx32 | multm_reduce_add3b0_maj3b_wy32;
  assign multm_reduce_add3b0_maj3b_or3b_wx33 = multm_reduce_add3b0_maj3b_wx33 | multm_reduce_add3b0_maj3b_wy33;
  assign multm_reduce_add3b0_maj3b_or3b_wx34 = multm_reduce_add3b0_maj3b_wx34 | multm_reduce_add3b0_maj3b_wy34;
  assign multm_reduce_add3b0_maj3b_or3b_wx35 = multm_reduce_add3b0_maj3b_wx35 | multm_reduce_add3b0_maj3b_wy35;
  assign multm_reduce_add3b0_maj3b_or3b_wx36 = multm_reduce_add3b0_maj3b_wx36 | multm_reduce_add3b0_maj3b_wy36;
  assign multm_reduce_add3b0_maj3b_or3b_wx37 = multm_reduce_add3b0_maj3b_wx37 | multm_reduce_add3b0_maj3b_wy37;
  assign multm_reduce_add3b0_maj3b_or3b_wx38 = multm_reduce_add3b0_maj3b_wx38 | multm_reduce_add3b0_maj3b_wy38;
  assign multm_reduce_add3b0_maj3b_or3b_wx39 = multm_reduce_add3b0_maj3b_wx39 | multm_reduce_add3b0_maj3b_wy39;
  assign multm_reduce_add3b0_maj3b_or3b_wx40 = multm_reduce_add3b0_maj3b_wx40 | multm_reduce_add3b0_maj3b_wy40;
  assign multm_reduce_add3b0_maj3b_or3b_wx41 = multm_reduce_add3b0_maj3b_wx41 | multm_reduce_add3b0_maj3b_wy41;
  assign multm_reduce_add3b0_maj3b_or3b_wx42 = multm_reduce_add3b0_maj3b_wx42 | multm_reduce_add3b0_maj3b_wy42;
  assign multm_reduce_add3b0_maj3b_or3b_wx43 = multm_reduce_add3b0_maj3b_wx43 | multm_reduce_add3b0_maj3b_wy43;
  assign multm_reduce_add3b0_maj3b_or3b_wx44 = multm_reduce_add3b0_maj3b_wx44 | multm_reduce_add3b0_maj3b_wy44;
  assign multm_reduce_add3b0_maj3b_or3b_wx45 = multm_reduce_add3b0_maj3b_wx45 | multm_reduce_add3b0_maj3b_wy45;
  assign multm_reduce_add3b0_maj3b_or3b_wx46 = multm_reduce_add3b0_maj3b_wx46 | multm_reduce_add3b0_maj3b_wy46;
  assign multm_reduce_add3b0_maj3b_or3b_wx47 = multm_reduce_add3b0_maj3b_wx47 | multm_reduce_add3b0_maj3b_wy47;
  assign multm_reduce_add3b0_maj3b_or3b_wx48 = multm_reduce_add3b0_maj3b_wx48 | multm_reduce_add3b0_maj3b_wy48;
  assign multm_reduce_add3b0_maj3b_or3b_wx49 = multm_reduce_add3b0_maj3b_wx49 | multm_reduce_add3b0_maj3b_wy49;
  assign multm_reduce_add3b0_maj3b_or3b_wx50 = multm_reduce_add3b0_maj3b_wx50 | multm_reduce_add3b0_maj3b_wy50;
  assign multm_reduce_add3b0_maj3b_or3b_wx51 = multm_reduce_add3b0_maj3b_wx51 | multm_reduce_add3b0_maj3b_wy51;
  assign multm_reduce_add3b0_maj3b_or3b_wx52 = multm_reduce_add3b0_maj3b_wx52 | multm_reduce_add3b0_maj3b_wy52;
  assign multm_reduce_add3b0_maj3b_or3b_wx53 = multm_reduce_add3b0_maj3b_wx53 | multm_reduce_add3b0_maj3b_wy53;
  assign multm_reduce_add3b0_maj3b_or3b_wx54 = multm_reduce_add3b0_maj3b_wx54 | multm_reduce_add3b0_maj3b_wy54;
  assign multm_reduce_add3b0_maj3b_or3b_wx55 = multm_reduce_add3b0_maj3b_wx55 | multm_reduce_add3b0_maj3b_wy55;
  assign multm_reduce_add3b0_maj3b_or3b_wx56 = multm_reduce_add3b0_maj3b_wx56 | multm_reduce_add3b0_maj3b_wy56;
  assign multm_reduce_add3b0_maj3b_or3b_wx57 = multm_reduce_add3b0_maj3b_wx57 | multm_reduce_add3b0_maj3b_wy57;
  assign multm_reduce_add3b0_maj3b_or3b_wx58 = multm_reduce_add3b0_maj3b_wx58 | multm_reduce_add3b0_maj3b_wy58;
  assign multm_reduce_add3b0_maj3b_or3b_wx59 = multm_reduce_add3b0_maj3b_wx59 | multm_reduce_add3b0_maj3b_wy59;
  assign multm_reduce_add3b0_maj3b_or3b_wx60 = multm_reduce_add3b0_maj3b_wx60 | multm_reduce_add3b0_maj3b_wy60;
  assign multm_reduce_add3b0_maj3b_or3b_wx61 = multm_reduce_add3b0_maj3b_wx61 | multm_reduce_add3b0_maj3b_wy61;
  assign multm_reduce_add3b0_maj3b_or3b_wx62 = multm_reduce_add3b0_maj3b_wx62 | multm_reduce_add3b0_maj3b_wy62;
  assign multm_reduce_add3b0_maj3b_or3b_wx63 = multm_reduce_add3b0_maj3b_wx63 | multm_reduce_add3b0_maj3b_wy63;
  assign multm_reduce_add3b0_maj3b_or3b_wx64 = multm_reduce_add3b0_maj3b_wx64 | multm_reduce_add3b0_maj3b_wy64;
  assign multm_reduce_add3b0_maj3b_or3b_wx65 = multm_reduce_add3b0_maj3b_wx65 | multm_reduce_add3b0_maj3b_wy65;
  assign multm_reduce_add3b0_maj3b_or3b_wx66 = multm_reduce_add3b0_maj3b_wx66 | multm_reduce_add3b0_maj3b_wy66;
  assign multm_reduce_add3b0_maj3b_or3b_wx67 = multm_reduce_add3b0_maj3b_wx67 | multm_reduce_add3b0_maj3b_wy67;
  assign multm_reduce_add3b0_maj3b_or3b_wx68 = multm_reduce_add3b0_maj3b_wx68 | multm_reduce_add3b0_maj3b_wy68;
  assign multm_reduce_add3b0_maj3b_or3b_wx69 = multm_reduce_add3b0_maj3b_wx69 | multm_reduce_add3b0_maj3b_wy69;
  assign multm_reduce_add3b0_maj3b_or3b_wx70 = multm_reduce_add3b0_maj3b_wx70 | multm_reduce_add3b0_maj3b_wy70;
  assign multm_reduce_add3b0_maj3b_or3b_wx71 = multm_reduce_add3b0_maj3b_wx71 | multm_reduce_add3b0_maj3b_wy71;
  assign multm_reduce_add3b0_maj3b_or3b_wx72 = multm_reduce_add3b0_maj3b_wx72 | multm_reduce_add3b0_maj3b_wy72;
  assign multm_reduce_add3b0_maj3b_or3b_wx73 = multm_reduce_add3b0_maj3b_wx73 | multm_reduce_add3b0_maj3b_wy73;
  assign multm_reduce_add3b0_maj3b_or3b_wx74 = multm_reduce_add3b0_maj3b_wx74 | multm_reduce_add3b0_maj3b_wy74;
  assign multm_reduce_add3b0_maj3b_or3b_wx75 = multm_reduce_add3b0_maj3b_wx75 | multm_reduce_add3b0_maj3b_wy75;
  assign multm_reduce_add3b0_maj3b_or3b_wx76 = multm_reduce_add3b0_maj3b_wx76 | multm_reduce_add3b0_maj3b_wy76;
  assign multm_reduce_add3b0_maj3b_or3b_wx77 = multm_reduce_add3b0_maj3b_wx77 | multm_reduce_add3b0_maj3b_wy77;
  assign multm_reduce_add3b0_maj3b_or3b_wx78 = multm_reduce_add3b0_maj3b_wx78 | multm_reduce_add3b0_maj3b_wy78;
  assign multm_reduce_add3b0_maj3b_or3b_wx79 = multm_reduce_add3b0_maj3b_wx79 | multm_reduce_add3b0_maj3b_wy79;
  assign multm_reduce_add3b0_maj3b_or3b_wx80 = multm_reduce_add3b0_maj3b_wx80 | multm_reduce_add3b0_maj3b_wy80;
  assign multm_reduce_add3b0_maj3b_or3b_wx81 = multm_reduce_add3b0_maj3b_wx81 | multm_reduce_add3b0_maj3b_wy81;
  assign multm_reduce_add3b0_maj3b_or3b_wx82 = multm_reduce_add3b0_maj3b_wx82 | multm_reduce_add3b0_maj3b_wy82;
  assign multm_reduce_add3b0_maj3b_or3b_wx83 = multm_reduce_add3b0_maj3b_wx83 | multm_reduce_add3b0_maj3b_wy83;
  assign multm_reduce_add3b0_maj3b_or3b_wx84 = multm_reduce_add3b0_maj3b_wx84 | multm_reduce_add3b0_maj3b_wy84;
  assign multm_reduce_add3b0_maj3b_or3b_wx85 = multm_reduce_add3b0_maj3b_wx85 | multm_reduce_add3b0_maj3b_wy85;
  assign multm_reduce_add3b0_maj3b_or3b_wx86 = multm_reduce_add3b0_maj3b_wx86 | multm_reduce_add3b0_maj3b_wy86;
  assign multm_reduce_add3b0_maj3b_or3b_wx87 = multm_reduce_add3b0_maj3b_wx87 | multm_reduce_add3b0_maj3b_wy87;
  assign multm_reduce_add3b0_maj3b_or3b_wx88 = multm_reduce_add3b0_maj3b_wx88 | multm_reduce_add3b0_maj3b_wy88;
  assign multm_reduce_add3b0_maj3b_or3b_wx89 = multm_reduce_add3b0_maj3b_wx89 | multm_reduce_add3b0_maj3b_wy89;
  assign multm_reduce_add3b0_maj3b_or3b_wx90 = multm_reduce_add3b0_maj3b_wx90 | multm_reduce_add3b0_maj3b_wy90;
  assign multm_reduce_add3b0_maj3b_or3b_wx91 = multm_reduce_add3b0_maj3b_wx91 | multm_reduce_add3b0_maj3b_wy91;
  assign multm_reduce_add3b0_maj3b_or3b_wx92 = multm_reduce_add3b0_maj3b_wx92 | multm_reduce_add3b0_maj3b_wy92;
  assign multm_reduce_add3b0_maj3b_or3b_wx93 = multm_reduce_add3b0_maj3b_wx93 | multm_reduce_add3b0_maj3b_wy93;
  assign multm_reduce_add3b0_maj3b_or3b_wx94 = multm_reduce_add3b0_maj3b_wx94 | multm_reduce_add3b0_maj3b_wy94;
  assign multm_reduce_add3b0_maj3b_or3b_wx95 = multm_reduce_add3b0_maj3b_wx95 | multm_reduce_add3b0_maj3b_wy95;
  assign multm_reduce_add3b0_maj3b_or3b_wx96 = multm_reduce_add3b0_maj3b_wx96 | multm_reduce_add3b0_maj3b_wy96;
  assign multm_reduce_add3b0_maj3b_or3b_wx97 = multm_reduce_add3b0_maj3b_wx97 | multm_reduce_add3b0_maj3b_wy97;
  assign multm_reduce_add3b0_maj3b_or3b_wx98 = multm_reduce_add3b0_maj3b_wx98 | multm_reduce_add3b0_maj3b_wy98;
  assign multm_reduce_add3b0_maj3b_or3b_wx99 = multm_reduce_add3b0_maj3b_wx99 | multm_reduce_add3b0_maj3b_wy99;
  assign multm_reduce_add3b0_maj3b_or3b_wx100 = multm_reduce_add3b0_maj3b_wx100 | multm_reduce_add3b0_maj3b_wy100;
  assign multm_reduce_add3b0_maj3b_or3b_wx101 = multm_reduce_add3b0_maj3b_wx101 | multm_reduce_add3b0_maj3b_wy101;
  assign multm_reduce_add3b0_maj3b_or3b_wx102 = multm_reduce_add3b0_maj3b_wx102 | multm_reduce_add3b0_maj3b_wy102;
  assign multm_reduce_add3b0_maj3b_or3b_wx103 = multm_reduce_add3b0_maj3b_wx103 | multm_reduce_add3b0_maj3b_wy103;
  assign multm_reduce_add3b0_maj3b_or3b_wx104 = multm_reduce_add3b0_maj3b_wx104 | multm_reduce_add3b0_maj3b_wy104;
  assign multm_reduce_add3b0_maj3b_or3b_wx105 = multm_reduce_add3b0_maj3b_wx105 | multm_reduce_add3b0_maj3b_wy105;
  assign multm_reduce_add3b0_maj3b_or3b_wx106 = multm_reduce_add3b0_maj3b_wx106 | multm_reduce_add3b0_maj3b_wy106;
  assign multm_reduce_add3b0_maj3b_or3b_wx107 = multm_reduce_add3b0_maj3b_wx107 | multm_reduce_add3b0_maj3b_wy107;
  assign multm_reduce_add3b0_maj3b_or3b_wx108 = multm_reduce_add3b0_maj3b_wx108 | multm_reduce_add3b0_maj3b_wy108;
  assign multm_reduce_add3b0_maj3b_or3b_wx109 = multm_reduce_add3b0_maj3b_wx109 | multm_reduce_add3b0_maj3b_wy109;
  assign multm_reduce_add3b0_maj3b_or3b_wx110 = multm_reduce_add3b0_maj3b_wx110 | multm_reduce_add3b0_maj3b_wy110;
  assign multm_reduce_add3b0_maj3b_or3b_wx111 = multm_reduce_add3b0_maj3b_wx111 | multm_reduce_add3b0_maj3b_wy111;
  assign multm_reduce_add3b0_maj3b_or3b_wx112 = multm_reduce_add3b0_maj3b_wx112 | multm_reduce_add3b0_maj3b_wy112;
  assign multm_reduce_add3b0_maj3b_or3b_wx113 = multm_reduce_add3b0_maj3b_wx113 | multm_reduce_add3b0_maj3b_wy113;
  assign multm_reduce_add3b0_maj3b_or3b_wx114 = multm_reduce_add3b0_maj3b_wx114 | multm_reduce_add3b0_maj3b_wy114;
  assign multm_reduce_add3b0_maj3b_or3b_wx115 = multm_reduce_add3b0_maj3b_wx115 | multm_reduce_add3b0_maj3b_wy115;
  assign multm_reduce_add3b0_maj3b_or3b_wx116 = multm_reduce_add3b0_maj3b_wx116 | multm_reduce_add3b0_maj3b_wy116;
  assign multm_reduce_add3b0_maj3b_or3b_wx117 = multm_reduce_add3b0_maj3b_wx117 | multm_reduce_add3b0_maj3b_wy117;
  assign multm_reduce_add3b0_maj3b_or3b_wx118 = multm_reduce_add3b0_maj3b_wx118 | multm_reduce_add3b0_maj3b_wy118;
  assign multm_reduce_add3b0_maj3b_or3b_wx119 = multm_reduce_add3b0_maj3b_wx119 | multm_reduce_add3b0_maj3b_wy119;
  assign multm_reduce_add3b0_maj3b_or3b_wx120 = multm_reduce_add3b0_maj3b_wx120 | multm_reduce_add3b0_maj3b_wy120;
  assign multm_reduce_add3b0_maj3b_or3b_wx121 = multm_reduce_add3b0_maj3b_wx121 | multm_reduce_add3b0_maj3b_wy121;
  assign multm_reduce_add3b0_maj3b_or3b_wx122 = multm_reduce_add3b0_maj3b_wx122 | multm_reduce_add3b0_maj3b_wy122;
  assign multm_reduce_add3b0_maj3b_or3b_wx123 = multm_reduce_add3b0_maj3b_wx123 | multm_reduce_add3b0_maj3b_wy123;
  assign multm_reduce_add3b0_maj3b_or3b_wx124 = multm_reduce_add3b0_maj3b_wx124 | multm_reduce_add3b0_maj3b_wy124;
  assign multm_reduce_add3b0_maj3b_or3b_wx125 = multm_reduce_add3b0_maj3b_wx125 | multm_reduce_add3b0_maj3b_wy125;
  assign multm_reduce_add3b0_maj3b_or3b_wx126 = multm_reduce_add3b0_maj3b_wx126 | multm_reduce_add3b0_maj3b_wy126;
  assign multm_reduce_add3b0_maj3b_or3b_wx127 = multm_reduce_add3b0_maj3b_wx127 | multm_reduce_add3b0_maj3b_wy127;
  assign multm_reduce_add3b0_maj3b_or3b_wx128 = multm_reduce_add3b0_maj3b_wx128 | multm_reduce_add3b0_maj3b_wy128;
  assign multm_reduce_add3b0_maj3b_or3b_wx129 = multm_reduce_add3b0_maj3b_wx129 | multm_reduce_add3b0_maj3b_wy129;
  assign multm_reduce_add3b0_maj3b_or3b_wx130 = multm_reduce_add3b0_maj3b_wx130 | multm_reduce_add3b0_maj3b_wy130;
  assign multm_reduce_add3b0_maj3b_or3b_wx131 = multm_reduce_add3b0_maj3b_wx131 | multm_reduce_add3b0_maj3b_wy131;
  assign multm_reduce_add3b0_maj3b_or3b_wx132 = multm_reduce_add3b0_maj3b_wx132 | multm_reduce_add3b0_maj3b_wy132;
  assign multm_reduce_add3b0_maj3b_or3b_wx133 = multm_reduce_add3b0_maj3b_wx133 | multm_reduce_add3b0_maj3b_wy133;
  assign multm_reduce_add3b0_maj3b_or3b_wx134 = multm_reduce_add3b0_maj3b_wx134 | multm_reduce_add3b0_maj3b_wy134;
  assign multm_reduce_add3b0_maj3b_or3b_wx135 = multm_reduce_add3b0_maj3b_wx135 | multm_reduce_add3b0_maj3b_wy135;
  assign multm_reduce_add3b0_maj3b_or3b_wx136 = multm_reduce_add3b0_maj3b_wx136 | multm_reduce_add3b0_maj3b_wy136;
  assign multm_reduce_add3b0_maj3b_or3b_wx137 = multm_reduce_add3b0_maj3b_wx137 | multm_reduce_add3b0_maj3b_wy137;
  assign multm_reduce_add3b0_maj3b_or3b_wx138 = multm_reduce_add3b0_maj3b_wx138 | multm_reduce_add3b0_maj3b_wy138;
  assign multm_reduce_add3b0_maj3b_or3b_wx139 = multm_reduce_add3b0_maj3b_wx139 | multm_reduce_add3b0_maj3b_wy139;
  assign multm_reduce_add3b0_maj3b_or3b_wx140 = multm_reduce_add3b0_maj3b_wx140 | multm_reduce_add3b0_maj3b_wy140;
  assign multm_reduce_add3b0_maj3b_or3b_wx141 = multm_reduce_add3b0_maj3b_wx141 | multm_reduce_add3b0_maj3b_wy141;
  assign multm_reduce_add3b0_maj3b_or3b_wx142 = multm_reduce_add3b0_maj3b_wx142 | multm_reduce_add3b0_maj3b_wy142;
  assign multm_reduce_add3b0_maj3b_or3b_wx143 = multm_reduce_add3b0_maj3b_wx143 | multm_reduce_add3b0_maj3b_wy143;
  assign multm_reduce_add3b0_maj3b_or3b_wx144 = multm_reduce_add3b0_maj3b_wx144 | multm_reduce_add3b0_maj3b_wy144;
  assign multm_reduce_add3b0_maj3b_or3b_wx145 = multm_reduce_add3b0_maj3b_wx145 | multm_reduce_add3b0_maj3b_wy145;
  assign multm_reduce_add3b0_maj3b_or3b_wx146 = multm_reduce_add3b0_maj3b_wx146 | multm_reduce_add3b0_maj3b_wy146;
  assign multm_reduce_add3b0_maj3b_or3b_wx147 = multm_reduce_add3b0_maj3b_wx147 | multm_reduce_add3b0_maj3b_wy147;
  assign multm_reduce_add3b0_maj3b_or3b_wx148 = multm_reduce_add3b0_maj3b_wx148 | multm_reduce_add3b0_maj3b_wy148;
  assign multm_reduce_add3b0_maj3b_or3b_wx149 = multm_reduce_add3b0_maj3b_wx149 | multm_reduce_add3b0_maj3b_wy149;
  assign multm_reduce_add3b0_maj3b_or3b_wx150 = multm_reduce_add3b0_maj3b_wx150 | multm_reduce_add3b0_maj3b_wy150;
  assign multm_reduce_add3b0_maj3b_or3b_wx151 = multm_reduce_add3b0_maj3b_wx151 | multm_reduce_add3b0_maj3b_wy151;
  assign multm_reduce_add3b0_maj3b_or3b_wx152 = multm_reduce_add3b0_maj3b_wx152 | multm_reduce_add3b0_maj3b_wy152;
  assign multm_reduce_add3b0_maj3b_or3b_wx153 = multm_reduce_add3b0_maj3b_wx153 | multm_reduce_add3b0_maj3b_wy153;
  assign multm_reduce_add3b0_maj3b_or3b_wx154 = multm_reduce_add3b0_maj3b_wx154 | multm_reduce_add3b0_maj3b_wy154;
  assign multm_reduce_add3b0_maj3b_or3b_wx155 = multm_reduce_add3b0_maj3b_wx155 | multm_reduce_add3b0_maj3b_wy155;
  assign multm_reduce_add3b0_maj3b_or3b_wx156 = multm_reduce_add3b0_maj3b_wx156 | multm_reduce_add3b0_maj3b_wy156;
  assign multm_reduce_add3b0_maj3b_or3b_wx157 = multm_reduce_add3b0_maj3b_wx157 | multm_reduce_add3b0_maj3b_wy157;
  assign multm_reduce_add3b0_maj3b_or3b_wx158 = multm_reduce_add3b0_maj3b_wx158 | multm_reduce_add3b0_maj3b_wy158;
  assign multm_reduce_add3b0_maj3b_or3b_wx159 = multm_reduce_add3b0_maj3b_wx159 | multm_reduce_add3b0_maj3b_wy159;
  assign multm_reduce_add3b0_maj3b_or3b_wx160 = multm_reduce_add3b0_maj3b_wx160 | multm_reduce_add3b0_maj3b_wy160;
  assign multm_reduce_add3b0_maj3b_or3b_wx161 = multm_reduce_add3b0_maj3b_wx161 | multm_reduce_add3b0_maj3b_wy161;
  assign multm_reduce_add3b0_maj3b_or3b_wx162 = multm_reduce_add3b0_maj3b_wx162 | multm_reduce_add3b0_maj3b_wy162;
  assign multm_reduce_add3b0_maj3b_or3b_wx163 = multm_reduce_add3b0_maj3b_wx163 | multm_reduce_add3b0_maj3b_wy163;
  assign multm_reduce_add3b0_maj3b_or3b_wx164 = multm_reduce_add3b0_maj3b_wx164 | multm_reduce_add3b0_maj3b_wy164;
  assign multm_reduce_add3b0_maj3b_or3b_wx165 = multm_reduce_add3b0_maj3b_wx165 | multm_reduce_add3b0_maj3b_wy165;
  assign multm_reduce_add3b0_maj3b_or3b_wx166 = multm_reduce_add3b0_maj3b_wx166 | multm_reduce_add3b0_maj3b_wy166;
  assign multm_reduce_add3b0_maj3b_or3b_wx167 = multm_reduce_add3b0_maj3b_wx167 | multm_reduce_add3b0_maj3b_wy167;
  assign multm_reduce_add3b0_maj3b_or3b_wx168 = multm_reduce_add3b0_maj3b_wx168 | multm_reduce_add3b0_maj3b_wy168;
  assign multm_reduce_add3b0_maj3b_or3b_wx169 = multm_reduce_add3b0_maj3b_wx169 | multm_reduce_add3b0_maj3b_wy169;
  assign multm_reduce_add3b0_maj3b_or3b_wx170 = multm_reduce_add3b0_maj3b_wx170 | multm_reduce_add3b0_maj3b_wy170;
  assign multm_reduce_add3b0_maj3b_or3b_wx171 = multm_reduce_add3b0_maj3b_wx171 | multm_reduce_add3b0_maj3b_wy171;
  assign multm_reduce_add3b0_maj3b_or3b_wx172 = multm_reduce_add3b0_maj3b_wx172 | multm_reduce_add3b0_maj3b_wy172;
  assign multm_reduce_add3b0_maj3b_or3b_wx173 = multm_reduce_add3b0_maj3b_wx173 | multm_reduce_add3b0_maj3b_wy173;
  assign multm_reduce_add3b0_maj3b_or3b_wx174 = multm_reduce_add3b0_maj3b_wx174 | multm_reduce_add3b0_maj3b_wy174;
  assign multm_reduce_add3b0_maj3b_or3b_wx175 = multm_reduce_add3b0_maj3b_wx175 | multm_reduce_add3b0_maj3b_wy175;
  assign multm_reduce_add3b0_maj3b_or3b_wx176 = multm_reduce_add3b0_maj3b_wx176 | multm_reduce_add3b0_maj3b_wy176;
  assign multm_reduce_add3b0_maj3b_or3b_wx177 = multm_reduce_add3b0_maj3b_wx177 | multm_reduce_add3b0_maj3b_wy177;
  assign multm_reduce_add3b0_maj3b_or3b_wx178 = multm_reduce_add3b0_maj3b_wx178 | multm_reduce_add3b0_maj3b_wy178;
  assign multm_reduce_add3b0_maj3b_or3b_wx179 = multm_reduce_add3b0_maj3b_wx179 | multm_reduce_add3b0_maj3b_wy179;
  assign multm_reduce_add3b0_maj3b_or3b_wx180 = multm_reduce_add3b0_maj3b_wx180 | multm_reduce_add3b0_maj3b_wy180;
  assign multm_reduce_add3b0_maj3b_or3b_wx181 = multm_reduce_add3b0_maj3b_wx181 | multm_reduce_add3b0_maj3b_wy181;
  assign multm_reduce_add3b0_maj3b_or3b_wx182 = multm_reduce_add3b0_maj3b_wx182 | multm_reduce_add3b0_maj3b_wy182;
  assign multm_reduce_add3b0_maj3b_wx0 = multm_reduce_sa0 & multm_reduce_sc0;
  assign multm_reduce_add3b0_maj3b_wx1 = multm_reduce_sa1 & multm_reduce_sc1;
  assign multm_reduce_add3b0_maj3b_wx2 = multm_reduce_sa2 & multm_reduce_sc2;
  assign multm_reduce_add3b0_maj3b_wx3 = multm_reduce_sa3 & multm_reduce_sc3;
  assign multm_reduce_add3b0_maj3b_wx4 = multm_reduce_sa4 & multm_reduce_sc4;
  assign multm_reduce_add3b0_maj3b_wx5 = multm_reduce_sa5 & multm_reduce_sc5;
  assign multm_reduce_add3b0_maj3b_wx6 = multm_reduce_sa6 & multm_reduce_sc6;
  assign multm_reduce_add3b0_maj3b_wx7 = multm_reduce_sa7 & multm_reduce_sc7;
  assign multm_reduce_add3b0_maj3b_wx8 = multm_reduce_sa8 & multm_reduce_sc8;
  assign multm_reduce_add3b0_maj3b_wx9 = multm_reduce_sa9 & multm_reduce_sc9;
  assign multm_reduce_add3b0_maj3b_wx10 = multm_reduce_sa10 & multm_reduce_sc10;
  assign multm_reduce_add3b0_maj3b_wx11 = multm_reduce_sa11 & multm_reduce_sc11;
  assign multm_reduce_add3b0_maj3b_wx12 = multm_reduce_sa12 & multm_reduce_sc12;
  assign multm_reduce_add3b0_maj3b_wx13 = multm_reduce_sa13 & multm_reduce_sc13;
  assign multm_reduce_add3b0_maj3b_wx14 = multm_reduce_sa14 & multm_reduce_sc14;
  assign multm_reduce_add3b0_maj3b_wx15 = multm_reduce_sa15 & multm_reduce_sc15;
  assign multm_reduce_add3b0_maj3b_wx16 = multm_reduce_sa16 & multm_reduce_sc16;
  assign multm_reduce_add3b0_maj3b_wx17 = multm_reduce_sa17 & multm_reduce_sc17;
  assign multm_reduce_add3b0_maj3b_wx18 = multm_reduce_sa18 & multm_reduce_sc18;
  assign multm_reduce_add3b0_maj3b_wx19 = multm_reduce_sa19 & multm_reduce_sc19;
  assign multm_reduce_add3b0_maj3b_wx20 = multm_reduce_sa20 & multm_reduce_sc20;
  assign multm_reduce_add3b0_maj3b_wx21 = multm_reduce_sa21 & multm_reduce_sc21;
  assign multm_reduce_add3b0_maj3b_wx22 = multm_reduce_sa22 & multm_reduce_sc22;
  assign multm_reduce_add3b0_maj3b_wx23 = multm_reduce_sa23 & multm_reduce_sc23;
  assign multm_reduce_add3b0_maj3b_wx24 = multm_reduce_sa24 & multm_reduce_sc24;
  assign multm_reduce_add3b0_maj3b_wx25 = multm_reduce_sa25 & multm_reduce_sc25;
  assign multm_reduce_add3b0_maj3b_wx26 = multm_reduce_sa26 & multm_reduce_sc26;
  assign multm_reduce_add3b0_maj3b_wx27 = multm_reduce_sa27 & multm_reduce_sc27;
  assign multm_reduce_add3b0_maj3b_wx28 = multm_reduce_sa28 & multm_reduce_sc28;
  assign multm_reduce_add3b0_maj3b_wx29 = multm_reduce_sa29 & multm_reduce_sc29;
  assign multm_reduce_add3b0_maj3b_wx30 = multm_reduce_sa30 & multm_reduce_sc30;
  assign multm_reduce_add3b0_maj3b_wx31 = multm_reduce_sa31 & multm_reduce_sc31;
  assign multm_reduce_add3b0_maj3b_wx32 = multm_reduce_sa32 & multm_reduce_sc32;
  assign multm_reduce_add3b0_maj3b_wx33 = multm_reduce_sa33 & multm_reduce_sc33;
  assign multm_reduce_add3b0_maj3b_wx34 = multm_reduce_sa34 & multm_reduce_sc34;
  assign multm_reduce_add3b0_maj3b_wx35 = multm_reduce_sa35 & multm_reduce_sc35;
  assign multm_reduce_add3b0_maj3b_wx36 = multm_reduce_sa36 & multm_reduce_sc36;
  assign multm_reduce_add3b0_maj3b_wx37 = multm_reduce_sa37 & multm_reduce_sc37;
  assign multm_reduce_add3b0_maj3b_wx38 = multm_reduce_sa38 & multm_reduce_sc38;
  assign multm_reduce_add3b0_maj3b_wx39 = multm_reduce_sa39 & multm_reduce_sc39;
  assign multm_reduce_add3b0_maj3b_wx40 = multm_reduce_sa40 & multm_reduce_sc40;
  assign multm_reduce_add3b0_maj3b_wx41 = multm_reduce_sa41 & multm_reduce_sc41;
  assign multm_reduce_add3b0_maj3b_wx42 = multm_reduce_sa42 & multm_reduce_sc42;
  assign multm_reduce_add3b0_maj3b_wx43 = multm_reduce_sa43 & multm_reduce_sc43;
  assign multm_reduce_add3b0_maj3b_wx44 = multm_reduce_sa44 & multm_reduce_sc44;
  assign multm_reduce_add3b0_maj3b_wx45 = multm_reduce_sa45 & multm_reduce_sc45;
  assign multm_reduce_add3b0_maj3b_wx46 = multm_reduce_sa46 & multm_reduce_sc46;
  assign multm_reduce_add3b0_maj3b_wx47 = multm_reduce_sa47 & multm_reduce_sc47;
  assign multm_reduce_add3b0_maj3b_wx48 = multm_reduce_sa48 & multm_reduce_sc48;
  assign multm_reduce_add3b0_maj3b_wx49 = multm_reduce_sa49 & multm_reduce_sc49;
  assign multm_reduce_add3b0_maj3b_wx50 = multm_reduce_sa50 & multm_reduce_sc50;
  assign multm_reduce_add3b0_maj3b_wx51 = multm_reduce_sa51 & multm_reduce_sc51;
  assign multm_reduce_add3b0_maj3b_wx52 = multm_reduce_sa52 & multm_reduce_sc52;
  assign multm_reduce_add3b0_maj3b_wx53 = multm_reduce_sa53 & multm_reduce_sc53;
  assign multm_reduce_add3b0_maj3b_wx54 = multm_reduce_sa54 & multm_reduce_sc54;
  assign multm_reduce_add3b0_maj3b_wx55 = multm_reduce_sa55 & multm_reduce_sc55;
  assign multm_reduce_add3b0_maj3b_wx56 = multm_reduce_sa56 & multm_reduce_sc56;
  assign multm_reduce_add3b0_maj3b_wx57 = multm_reduce_sa57 & multm_reduce_sc57;
  assign multm_reduce_add3b0_maj3b_wx58 = multm_reduce_sa58 & multm_reduce_sc58;
  assign multm_reduce_add3b0_maj3b_wx59 = multm_reduce_sa59 & multm_reduce_sc59;
  assign multm_reduce_add3b0_maj3b_wx60 = multm_reduce_sa60 & multm_reduce_sc60;
  assign multm_reduce_add3b0_maj3b_wx61 = multm_reduce_sa61 & multm_reduce_sc61;
  assign multm_reduce_add3b0_maj3b_wx62 = multm_reduce_sa62 & multm_reduce_sc62;
  assign multm_reduce_add3b0_maj3b_wx63 = multm_reduce_sa63 & multm_reduce_sc63;
  assign multm_reduce_add3b0_maj3b_wx64 = multm_reduce_sa64 & multm_reduce_sc64;
  assign multm_reduce_add3b0_maj3b_wx65 = multm_reduce_sa65 & multm_reduce_sc65;
  assign multm_reduce_add3b0_maj3b_wx66 = multm_reduce_sa66 & multm_reduce_sc66;
  assign multm_reduce_add3b0_maj3b_wx67 = multm_reduce_sa67 & multm_reduce_sc67;
  assign multm_reduce_add3b0_maj3b_wx68 = multm_reduce_sa68 & multm_reduce_sc68;
  assign multm_reduce_add3b0_maj3b_wx69 = multm_reduce_sa69 & multm_reduce_sc69;
  assign multm_reduce_add3b0_maj3b_wx70 = multm_reduce_sa70 & multm_reduce_sc70;
  assign multm_reduce_add3b0_maj3b_wx71 = multm_reduce_sa71 & multm_reduce_sc71;
  assign multm_reduce_add3b0_maj3b_wx72 = multm_reduce_sa72 & multm_reduce_sc72;
  assign multm_reduce_add3b0_maj3b_wx73 = multm_reduce_sa73 & multm_reduce_sc73;
  assign multm_reduce_add3b0_maj3b_wx74 = multm_reduce_sa74 & multm_reduce_sc74;
  assign multm_reduce_add3b0_maj3b_wx75 = multm_reduce_sa75 & multm_reduce_sc75;
  assign multm_reduce_add3b0_maj3b_wx76 = multm_reduce_sa76 & multm_reduce_sc76;
  assign multm_reduce_add3b0_maj3b_wx77 = multm_reduce_sa77 & multm_reduce_sc77;
  assign multm_reduce_add3b0_maj3b_wx78 = multm_reduce_sa78 & multm_reduce_sc78;
  assign multm_reduce_add3b0_maj3b_wx79 = multm_reduce_sa79 & multm_reduce_sc79;
  assign multm_reduce_add3b0_maj3b_wx80 = multm_reduce_sa80 & multm_reduce_sc80;
  assign multm_reduce_add3b0_maj3b_wx81 = multm_reduce_sa81 & multm_reduce_sc81;
  assign multm_reduce_add3b0_maj3b_wx82 = multm_reduce_sa82 & multm_reduce_sc82;
  assign multm_reduce_add3b0_maj3b_wx83 = multm_reduce_sa83 & multm_reduce_sc83;
  assign multm_reduce_add3b0_maj3b_wx84 = multm_reduce_sa84 & multm_reduce_sc84;
  assign multm_reduce_add3b0_maj3b_wx85 = multm_reduce_sa85 & multm_reduce_sc85;
  assign multm_reduce_add3b0_maj3b_wx86 = multm_reduce_sa86 & multm_reduce_sc86;
  assign multm_reduce_add3b0_maj3b_wx87 = multm_reduce_sa87 & multm_reduce_sc87;
  assign multm_reduce_add3b0_maj3b_wx88 = multm_reduce_sa88 & multm_reduce_sc88;
  assign multm_reduce_add3b0_maj3b_wx89 = multm_reduce_sa89 & multm_reduce_sc89;
  assign multm_reduce_add3b0_maj3b_wx90 = multm_reduce_sa90 & multm_reduce_sc90;
  assign multm_reduce_add3b0_maj3b_wx91 = multm_reduce_sa91 & multm_reduce_sc91;
  assign multm_reduce_add3b0_maj3b_wx92 = multm_reduce_sa92 & multm_reduce_sc92;
  assign multm_reduce_add3b0_maj3b_wx93 = multm_reduce_sa93 & multm_reduce_sc93;
  assign multm_reduce_add3b0_maj3b_wx94 = multm_reduce_sa94 & multm_reduce_sc94;
  assign multm_reduce_add3b0_maj3b_wx95 = multm_reduce_sa95 & multm_reduce_sc95;
  assign multm_reduce_add3b0_maj3b_wx96 = multm_reduce_sa96 & multm_reduce_sc96;
  assign multm_reduce_add3b0_maj3b_wx97 = multm_reduce_sa97 & multm_reduce_sc97;
  assign multm_reduce_add3b0_maj3b_wx98 = multm_reduce_sa98 & multm_reduce_sc98;
  assign multm_reduce_add3b0_maj3b_wx99 = multm_reduce_sa99 & multm_reduce_sc99;
  assign multm_reduce_add3b0_maj3b_wx100 = multm_reduce_sa100 & multm_reduce_sc100;
  assign multm_reduce_add3b0_maj3b_wx101 = multm_reduce_sa101 & multm_reduce_sc101;
  assign multm_reduce_add3b0_maj3b_wx102 = multm_reduce_sa102 & multm_reduce_sc102;
  assign multm_reduce_add3b0_maj3b_wx103 = multm_reduce_sa103 & multm_reduce_sc103;
  assign multm_reduce_add3b0_maj3b_wx104 = multm_reduce_sa104 & multm_reduce_sc104;
  assign multm_reduce_add3b0_maj3b_wx105 = multm_reduce_sa105 & multm_reduce_sc105;
  assign multm_reduce_add3b0_maj3b_wx106 = multm_reduce_sa106 & multm_reduce_sc106;
  assign multm_reduce_add3b0_maj3b_wx107 = multm_reduce_sa107 & multm_reduce_sc107;
  assign multm_reduce_add3b0_maj3b_wx108 = multm_reduce_sa108 & multm_reduce_sc108;
  assign multm_reduce_add3b0_maj3b_wx109 = multm_reduce_sa109 & multm_reduce_sc109;
  assign multm_reduce_add3b0_maj3b_wx110 = multm_reduce_sa110 & multm_reduce_sc110;
  assign multm_reduce_add3b0_maj3b_wx111 = multm_reduce_sa111 & multm_reduce_sc111;
  assign multm_reduce_add3b0_maj3b_wx112 = multm_reduce_sa112 & multm_reduce_sc112;
  assign multm_reduce_add3b0_maj3b_wx113 = multm_reduce_sa113 & multm_reduce_sc113;
  assign multm_reduce_add3b0_maj3b_wx114 = multm_reduce_sa114 & multm_reduce_sc114;
  assign multm_reduce_add3b0_maj3b_wx115 = multm_reduce_sa115 & multm_reduce_sc115;
  assign multm_reduce_add3b0_maj3b_wx116 = multm_reduce_sa116 & multm_reduce_sc116;
  assign multm_reduce_add3b0_maj3b_wx117 = multm_reduce_sa117 & multm_reduce_sc117;
  assign multm_reduce_add3b0_maj3b_wx118 = multm_reduce_sa118 & multm_reduce_sc118;
  assign multm_reduce_add3b0_maj3b_wx119 = multm_reduce_sa119 & multm_reduce_sc119;
  assign multm_reduce_add3b0_maj3b_wx120 = multm_reduce_sa120 & multm_reduce_sc120;
  assign multm_reduce_add3b0_maj3b_wx121 = multm_reduce_sa121 & multm_reduce_sc121;
  assign multm_reduce_add3b0_maj3b_wx122 = multm_reduce_sa122 & multm_reduce_sc122;
  assign multm_reduce_add3b0_maj3b_wx123 = multm_reduce_sa123 & multm_reduce_sc123;
  assign multm_reduce_add3b0_maj3b_wx124 = multm_reduce_sa124 & multm_reduce_sc124;
  assign multm_reduce_add3b0_maj3b_wx125 = multm_reduce_sa125 & multm_reduce_sc125;
  assign multm_reduce_add3b0_maj3b_wx126 = multm_reduce_sa126 & multm_reduce_sc126;
  assign multm_reduce_add3b0_maj3b_wx127 = multm_reduce_sa127 & multm_reduce_sc127;
  assign multm_reduce_add3b0_maj3b_wx128 = multm_reduce_sa128 & multm_reduce_sc128;
  assign multm_reduce_add3b0_maj3b_wx129 = multm_reduce_sa129 & multm_reduce_sc129;
  assign multm_reduce_add3b0_maj3b_wx130 = multm_reduce_sa130 & multm_reduce_sc130;
  assign multm_reduce_add3b0_maj3b_wx131 = multm_reduce_sa131 & multm_reduce_sc131;
  assign multm_reduce_add3b0_maj3b_wx132 = multm_reduce_sa132 & multm_reduce_sc132;
  assign multm_reduce_add3b0_maj3b_wx133 = multm_reduce_sa133 & multm_reduce_sc133;
  assign multm_reduce_add3b0_maj3b_wx134 = multm_reduce_sa134 & multm_reduce_sc134;
  assign multm_reduce_add3b0_maj3b_wx135 = multm_reduce_sa135 & multm_reduce_sc135;
  assign multm_reduce_add3b0_maj3b_wx136 = multm_reduce_sa136 & multm_reduce_sc136;
  assign multm_reduce_add3b0_maj3b_wx137 = multm_reduce_sa137 & multm_reduce_sc137;
  assign multm_reduce_add3b0_maj3b_wx138 = multm_reduce_sa138 & multm_reduce_sc138;
  assign multm_reduce_add3b0_maj3b_wx139 = multm_reduce_sa139 & multm_reduce_sc139;
  assign multm_reduce_add3b0_maj3b_wx140 = multm_reduce_sa140 & multm_reduce_sc140;
  assign multm_reduce_add3b0_maj3b_wx141 = multm_reduce_sa141 & multm_reduce_sc141;
  assign multm_reduce_add3b0_maj3b_wx142 = multm_reduce_sa142 & multm_reduce_sc142;
  assign multm_reduce_add3b0_maj3b_wx143 = multm_reduce_sa143 & multm_reduce_sc143;
  assign multm_reduce_add3b0_maj3b_wx144 = multm_reduce_sa144 & multm_reduce_sc144;
  assign multm_reduce_add3b0_maj3b_wx145 = multm_reduce_sa145 & multm_reduce_sc145;
  assign multm_reduce_add3b0_maj3b_wx146 = multm_reduce_sa146 & multm_reduce_sc146;
  assign multm_reduce_add3b0_maj3b_wx147 = multm_reduce_sa147 & multm_reduce_sc147;
  assign multm_reduce_add3b0_maj3b_wx148 = multm_reduce_sa148 & multm_reduce_sc148;
  assign multm_reduce_add3b0_maj3b_wx149 = multm_reduce_sa149 & multm_reduce_sc149;
  assign multm_reduce_add3b0_maj3b_wx150 = multm_reduce_sa150 & multm_reduce_sc150;
  assign multm_reduce_add3b0_maj3b_wx151 = multm_reduce_sa151 & multm_reduce_sc151;
  assign multm_reduce_add3b0_maj3b_wx152 = multm_reduce_sa152 & multm_reduce_sc152;
  assign multm_reduce_add3b0_maj3b_wx153 = multm_reduce_sa153 & multm_reduce_sc153;
  assign multm_reduce_add3b0_maj3b_wx154 = multm_reduce_sa154 & multm_reduce_sc154;
  assign multm_reduce_add3b0_maj3b_wx155 = multm_reduce_sa155 & multm_reduce_sc155;
  assign multm_reduce_add3b0_maj3b_wx156 = multm_reduce_sa156 & multm_reduce_sc156;
  assign multm_reduce_add3b0_maj3b_wx157 = multm_reduce_sa157 & multm_reduce_sc157;
  assign multm_reduce_add3b0_maj3b_wx158 = multm_reduce_sa158 & multm_reduce_sc158;
  assign multm_reduce_add3b0_maj3b_wx159 = multm_reduce_sa159 & multm_reduce_sc159;
  assign multm_reduce_add3b0_maj3b_wx160 = multm_reduce_sa160 & multm_reduce_sc160;
  assign multm_reduce_add3b0_maj3b_wx161 = multm_reduce_sa161 & multm_reduce_sc161;
  assign multm_reduce_add3b0_maj3b_wx162 = multm_reduce_sa162 & multm_reduce_sc162;
  assign multm_reduce_add3b0_maj3b_wx163 = multm_reduce_sa163 & multm_reduce_sc163;
  assign multm_reduce_add3b0_maj3b_wx164 = multm_reduce_sa164 & multm_reduce_sc164;
  assign multm_reduce_add3b0_maj3b_wx165 = multm_reduce_sa165 & multm_reduce_sc165;
  assign multm_reduce_add3b0_maj3b_wx166 = multm_reduce_sa166 & multm_reduce_sc166;
  assign multm_reduce_add3b0_maj3b_wx167 = multm_reduce_sa167 & multm_reduce_sc167;
  assign multm_reduce_add3b0_maj3b_wx168 = multm_reduce_sa168 & multm_reduce_sc168;
  assign multm_reduce_add3b0_maj3b_wx169 = multm_reduce_sa169 & multm_reduce_sc169;
  assign multm_reduce_add3b0_maj3b_wx170 = multm_reduce_sa170 & multm_reduce_sc170;
  assign multm_reduce_add3b0_maj3b_wx171 = multm_reduce_sa171 & multm_reduce_sc171;
  assign multm_reduce_add3b0_maj3b_wx172 = multm_reduce_sa172 & multm_reduce_sc172;
  assign multm_reduce_add3b0_maj3b_wx173 = multm_reduce_sa173 & multm_reduce_sc173;
  assign multm_reduce_add3b0_maj3b_wx174 = multm_reduce_sa174 & multm_reduce_sc174;
  assign multm_reduce_add3b0_maj3b_wx175 = multm_reduce_sa175 & multm_reduce_sc175;
  assign multm_reduce_add3b0_maj3b_wx176 = multm_reduce_sa176 & multm_reduce_sc176;
  assign multm_reduce_add3b0_maj3b_wx177 = multm_reduce_sa177 & multm_reduce_sc177;
  assign multm_reduce_add3b0_maj3b_wx178 = multm_reduce_sa178 & multm_reduce_sc178;
  assign multm_reduce_add3b0_maj3b_wx179 = multm_reduce_sa179 & multm_reduce_sc179;
  assign multm_reduce_add3b0_maj3b_wx180 = multm_reduce_sa180 & multm_reduce_sc180;
  assign multm_reduce_add3b0_maj3b_wx181 = multm_reduce_sa181 & multm_reduce_sc181;
  assign multm_reduce_add3b0_maj3b_wx182 = multm_reduce_sa182 & multm_reduce_sc182;
  assign multm_reduce_add3b0_maj3b_wy0 = multm_reduce_sa0 & multm_reduce_sd0;
  assign multm_reduce_add3b0_maj3b_wy1 = multm_reduce_sa1 & multm_reduce_sd1;
  assign multm_reduce_add3b0_maj3b_wy2 = multm_reduce_sa2 & multm_reduce_sd2;
  assign multm_reduce_add3b0_maj3b_wy3 = multm_reduce_sa3 & multm_reduce_sd3;
  assign multm_reduce_add3b0_maj3b_wy4 = multm_reduce_sa4 & multm_reduce_sd4;
  assign multm_reduce_add3b0_maj3b_wy5 = multm_reduce_sa5 & multm_reduce_sd5;
  assign multm_reduce_add3b0_maj3b_wy6 = multm_reduce_sa6 & multm_reduce_sd6;
  assign multm_reduce_add3b0_maj3b_wy7 = multm_reduce_sa7 & multm_reduce_sd7;
  assign multm_reduce_add3b0_maj3b_wy8 = multm_reduce_sa8 & multm_reduce_sd8;
  assign multm_reduce_add3b0_maj3b_wy9 = multm_reduce_sa9 & multm_reduce_sd9;
  assign multm_reduce_add3b0_maj3b_wy10 = multm_reduce_sa10 & multm_reduce_sd10;
  assign multm_reduce_add3b0_maj3b_wy11 = multm_reduce_sa11 & multm_reduce_sd11;
  assign multm_reduce_add3b0_maj3b_wy12 = multm_reduce_sa12 & multm_reduce_sd12;
  assign multm_reduce_add3b0_maj3b_wy13 = multm_reduce_sa13 & multm_reduce_sd13;
  assign multm_reduce_add3b0_maj3b_wy14 = multm_reduce_sa14 & multm_reduce_sd14;
  assign multm_reduce_add3b0_maj3b_wy15 = multm_reduce_sa15 & multm_reduce_sd15;
  assign multm_reduce_add3b0_maj3b_wy16 = multm_reduce_sa16 & multm_reduce_sd16;
  assign multm_reduce_add3b0_maj3b_wy17 = multm_reduce_sa17 & multm_reduce_sd17;
  assign multm_reduce_add3b0_maj3b_wy18 = multm_reduce_sa18 & multm_reduce_sd18;
  assign multm_reduce_add3b0_maj3b_wy19 = multm_reduce_sa19 & multm_reduce_sd19;
  assign multm_reduce_add3b0_maj3b_wy20 = multm_reduce_sa20 & multm_reduce_sd20;
  assign multm_reduce_add3b0_maj3b_wy21 = multm_reduce_sa21 & multm_reduce_sd21;
  assign multm_reduce_add3b0_maj3b_wy22 = multm_reduce_sa22 & multm_reduce_sd22;
  assign multm_reduce_add3b0_maj3b_wy23 = multm_reduce_sa23 & multm_reduce_sd23;
  assign multm_reduce_add3b0_maj3b_wy24 = multm_reduce_sa24 & multm_reduce_sd24;
  assign multm_reduce_add3b0_maj3b_wy25 = multm_reduce_sa25 & multm_reduce_sd25;
  assign multm_reduce_add3b0_maj3b_wy26 = multm_reduce_sa26 & multm_reduce_sd26;
  assign multm_reduce_add3b0_maj3b_wy27 = multm_reduce_sa27 & multm_reduce_sd27;
  assign multm_reduce_add3b0_maj3b_wy28 = multm_reduce_sa28 & multm_reduce_sd28;
  assign multm_reduce_add3b0_maj3b_wy29 = multm_reduce_sa29 & multm_reduce_sd29;
  assign multm_reduce_add3b0_maj3b_wy30 = multm_reduce_sa30 & multm_reduce_sd30;
  assign multm_reduce_add3b0_maj3b_wy31 = multm_reduce_sa31 & multm_reduce_sd31;
  assign multm_reduce_add3b0_maj3b_wy32 = multm_reduce_sa32 & multm_reduce_sd32;
  assign multm_reduce_add3b0_maj3b_wy33 = multm_reduce_sa33 & multm_reduce_sd33;
  assign multm_reduce_add3b0_maj3b_wy34 = multm_reduce_sa34 & multm_reduce_sd34;
  assign multm_reduce_add3b0_maj3b_wy35 = multm_reduce_sa35 & multm_reduce_sd35;
  assign multm_reduce_add3b0_maj3b_wy36 = multm_reduce_sa36 & multm_reduce_sd36;
  assign multm_reduce_add3b0_maj3b_wy37 = multm_reduce_sa37 & multm_reduce_sd37;
  assign multm_reduce_add3b0_maj3b_wy38 = multm_reduce_sa38 & multm_reduce_sd38;
  assign multm_reduce_add3b0_maj3b_wy39 = multm_reduce_sa39 & multm_reduce_sd39;
  assign multm_reduce_add3b0_maj3b_wy40 = multm_reduce_sa40 & multm_reduce_sd40;
  assign multm_reduce_add3b0_maj3b_wy41 = multm_reduce_sa41 & multm_reduce_sd41;
  assign multm_reduce_add3b0_maj3b_wy42 = multm_reduce_sa42 & multm_reduce_sd42;
  assign multm_reduce_add3b0_maj3b_wy43 = multm_reduce_sa43 & multm_reduce_sd43;
  assign multm_reduce_add3b0_maj3b_wy44 = multm_reduce_sa44 & multm_reduce_sd44;
  assign multm_reduce_add3b0_maj3b_wy45 = multm_reduce_sa45 & multm_reduce_sd45;
  assign multm_reduce_add3b0_maj3b_wy46 = multm_reduce_sa46 & multm_reduce_sd46;
  assign multm_reduce_add3b0_maj3b_wy47 = multm_reduce_sa47 & multm_reduce_sd47;
  assign multm_reduce_add3b0_maj3b_wy48 = multm_reduce_sa48 & multm_reduce_sd48;
  assign multm_reduce_add3b0_maj3b_wy49 = multm_reduce_sa49 & multm_reduce_sd49;
  assign multm_reduce_add3b0_maj3b_wy50 = multm_reduce_sa50 & multm_reduce_sd50;
  assign multm_reduce_add3b0_maj3b_wy51 = multm_reduce_sa51 & multm_reduce_sd51;
  assign multm_reduce_add3b0_maj3b_wy52 = multm_reduce_sa52 & multm_reduce_sd52;
  assign multm_reduce_add3b0_maj3b_wy53 = multm_reduce_sa53 & multm_reduce_sd53;
  assign multm_reduce_add3b0_maj3b_wy54 = multm_reduce_sa54 & multm_reduce_sd54;
  assign multm_reduce_add3b0_maj3b_wy55 = multm_reduce_sa55 & multm_reduce_sd55;
  assign multm_reduce_add3b0_maj3b_wy56 = multm_reduce_sa56 & multm_reduce_sd56;
  assign multm_reduce_add3b0_maj3b_wy57 = multm_reduce_sa57 & multm_reduce_sd57;
  assign multm_reduce_add3b0_maj3b_wy58 = multm_reduce_sa58 & multm_reduce_sd58;
  assign multm_reduce_add3b0_maj3b_wy59 = multm_reduce_sa59 & multm_reduce_sd59;
  assign multm_reduce_add3b0_maj3b_wy60 = multm_reduce_sa60 & multm_reduce_sd60;
  assign multm_reduce_add3b0_maj3b_wy61 = multm_reduce_sa61 & multm_reduce_sd61;
  assign multm_reduce_add3b0_maj3b_wy62 = multm_reduce_sa62 & multm_reduce_sd62;
  assign multm_reduce_add3b0_maj3b_wy63 = multm_reduce_sa63 & multm_reduce_sd63;
  assign multm_reduce_add3b0_maj3b_wy64 = multm_reduce_sa64 & multm_reduce_sd64;
  assign multm_reduce_add3b0_maj3b_wy65 = multm_reduce_sa65 & multm_reduce_sd65;
  assign multm_reduce_add3b0_maj3b_wy66 = multm_reduce_sa66 & multm_reduce_sd66;
  assign multm_reduce_add3b0_maj3b_wy67 = multm_reduce_sa67 & multm_reduce_sd67;
  assign multm_reduce_add3b0_maj3b_wy68 = multm_reduce_sa68 & multm_reduce_sd68;
  assign multm_reduce_add3b0_maj3b_wy69 = multm_reduce_sa69 & multm_reduce_sd69;
  assign multm_reduce_add3b0_maj3b_wy70 = multm_reduce_sa70 & multm_reduce_sd70;
  assign multm_reduce_add3b0_maj3b_wy71 = multm_reduce_sa71 & multm_reduce_sd71;
  assign multm_reduce_add3b0_maj3b_wy72 = multm_reduce_sa72 & multm_reduce_sd72;
  assign multm_reduce_add3b0_maj3b_wy73 = multm_reduce_sa73 & multm_reduce_sd73;
  assign multm_reduce_add3b0_maj3b_wy74 = multm_reduce_sa74 & multm_reduce_sd74;
  assign multm_reduce_add3b0_maj3b_wy75 = multm_reduce_sa75 & multm_reduce_sd75;
  assign multm_reduce_add3b0_maj3b_wy76 = multm_reduce_sa76 & multm_reduce_sd76;
  assign multm_reduce_add3b0_maj3b_wy77 = multm_reduce_sa77 & multm_reduce_sd77;
  assign multm_reduce_add3b0_maj3b_wy78 = multm_reduce_sa78 & multm_reduce_sd78;
  assign multm_reduce_add3b0_maj3b_wy79 = multm_reduce_sa79 & multm_reduce_sd79;
  assign multm_reduce_add3b0_maj3b_wy80 = multm_reduce_sa80 & multm_reduce_sd80;
  assign multm_reduce_add3b0_maj3b_wy81 = multm_reduce_sa81 & multm_reduce_sd81;
  assign multm_reduce_add3b0_maj3b_wy82 = multm_reduce_sa82 & multm_reduce_sd82;
  assign multm_reduce_add3b0_maj3b_wy83 = multm_reduce_sa83 & multm_reduce_sd83;
  assign multm_reduce_add3b0_maj3b_wy84 = multm_reduce_sa84 & multm_reduce_sd84;
  assign multm_reduce_add3b0_maj3b_wy85 = multm_reduce_sa85 & multm_reduce_sd85;
  assign multm_reduce_add3b0_maj3b_wy86 = multm_reduce_sa86 & multm_reduce_sd86;
  assign multm_reduce_add3b0_maj3b_wy87 = multm_reduce_sa87 & multm_reduce_sd87;
  assign multm_reduce_add3b0_maj3b_wy88 = multm_reduce_sa88 & multm_reduce_sd88;
  assign multm_reduce_add3b0_maj3b_wy89 = multm_reduce_sa89 & multm_reduce_sd89;
  assign multm_reduce_add3b0_maj3b_wy90 = multm_reduce_sa90 & multm_reduce_sd90;
  assign multm_reduce_add3b0_maj3b_wy91 = multm_reduce_sa91 & multm_reduce_sd91;
  assign multm_reduce_add3b0_maj3b_wy92 = multm_reduce_sa92 & multm_reduce_sd92;
  assign multm_reduce_add3b0_maj3b_wy93 = multm_reduce_sa93 & multm_reduce_sd93;
  assign multm_reduce_add3b0_maj3b_wy94 = multm_reduce_sa94 & multm_reduce_sd94;
  assign multm_reduce_add3b0_maj3b_wy95 = multm_reduce_sa95 & multm_reduce_sd95;
  assign multm_reduce_add3b0_maj3b_wy96 = multm_reduce_sa96 & multm_reduce_sd96;
  assign multm_reduce_add3b0_maj3b_wy97 = multm_reduce_sa97 & multm_reduce_sd97;
  assign multm_reduce_add3b0_maj3b_wy98 = multm_reduce_sa98 & multm_reduce_sd98;
  assign multm_reduce_add3b0_maj3b_wy99 = multm_reduce_sa99 & multm_reduce_sd99;
  assign multm_reduce_add3b0_maj3b_wy100 = multm_reduce_sa100 & multm_reduce_sd100;
  assign multm_reduce_add3b0_maj3b_wy101 = multm_reduce_sa101 & multm_reduce_sd101;
  assign multm_reduce_add3b0_maj3b_wy102 = multm_reduce_sa102 & multm_reduce_sd102;
  assign multm_reduce_add3b0_maj3b_wy103 = multm_reduce_sa103 & multm_reduce_sd103;
  assign multm_reduce_add3b0_maj3b_wy104 = multm_reduce_sa104 & multm_reduce_sd104;
  assign multm_reduce_add3b0_maj3b_wy105 = multm_reduce_sa105 & multm_reduce_sd105;
  assign multm_reduce_add3b0_maj3b_wy106 = multm_reduce_sa106 & multm_reduce_sd106;
  assign multm_reduce_add3b0_maj3b_wy107 = multm_reduce_sa107 & multm_reduce_sd107;
  assign multm_reduce_add3b0_maj3b_wy108 = multm_reduce_sa108 & multm_reduce_sd108;
  assign multm_reduce_add3b0_maj3b_wy109 = multm_reduce_sa109 & multm_reduce_sd109;
  assign multm_reduce_add3b0_maj3b_wy110 = multm_reduce_sa110 & multm_reduce_sd110;
  assign multm_reduce_add3b0_maj3b_wy111 = multm_reduce_sa111 & multm_reduce_sd111;
  assign multm_reduce_add3b0_maj3b_wy112 = multm_reduce_sa112 & multm_reduce_sd112;
  assign multm_reduce_add3b0_maj3b_wy113 = multm_reduce_sa113 & multm_reduce_sd113;
  assign multm_reduce_add3b0_maj3b_wy114 = multm_reduce_sa114 & multm_reduce_sd114;
  assign multm_reduce_add3b0_maj3b_wy115 = multm_reduce_sa115 & multm_reduce_sd115;
  assign multm_reduce_add3b0_maj3b_wy116 = multm_reduce_sa116 & multm_reduce_sd116;
  assign multm_reduce_add3b0_maj3b_wy117 = multm_reduce_sa117 & multm_reduce_sd117;
  assign multm_reduce_add3b0_maj3b_wy118 = multm_reduce_sa118 & multm_reduce_sd118;
  assign multm_reduce_add3b0_maj3b_wy119 = multm_reduce_sa119 & multm_reduce_sd119;
  assign multm_reduce_add3b0_maj3b_wy120 = multm_reduce_sa120 & multm_reduce_sd120;
  assign multm_reduce_add3b0_maj3b_wy121 = multm_reduce_sa121 & multm_reduce_sd121;
  assign multm_reduce_add3b0_maj3b_wy122 = multm_reduce_sa122 & multm_reduce_sd122;
  assign multm_reduce_add3b0_maj3b_wy123 = multm_reduce_sa123 & multm_reduce_sd123;
  assign multm_reduce_add3b0_maj3b_wy124 = multm_reduce_sa124 & multm_reduce_sd124;
  assign multm_reduce_add3b0_maj3b_wy125 = multm_reduce_sa125 & multm_reduce_sd125;
  assign multm_reduce_add3b0_maj3b_wy126 = multm_reduce_sa126 & multm_reduce_sd126;
  assign multm_reduce_add3b0_maj3b_wy127 = multm_reduce_sa127 & multm_reduce_sd127;
  assign multm_reduce_add3b0_maj3b_wy128 = multm_reduce_sa128 & multm_reduce_sd128;
  assign multm_reduce_add3b0_maj3b_wy129 = multm_reduce_sa129 & multm_reduce_sd129;
  assign multm_reduce_add3b0_maj3b_wy130 = multm_reduce_sa130 & multm_reduce_sd130;
  assign multm_reduce_add3b0_maj3b_wy131 = multm_reduce_sa131 & multm_reduce_sd131;
  assign multm_reduce_add3b0_maj3b_wy132 = multm_reduce_sa132 & multm_reduce_sd132;
  assign multm_reduce_add3b0_maj3b_wy133 = multm_reduce_sa133 & multm_reduce_sd133;
  assign multm_reduce_add3b0_maj3b_wy134 = multm_reduce_sa134 & multm_reduce_sd134;
  assign multm_reduce_add3b0_maj3b_wy135 = multm_reduce_sa135 & multm_reduce_sd135;
  assign multm_reduce_add3b0_maj3b_wy136 = multm_reduce_sa136 & multm_reduce_sd136;
  assign multm_reduce_add3b0_maj3b_wy137 = multm_reduce_sa137 & multm_reduce_sd137;
  assign multm_reduce_add3b0_maj3b_wy138 = multm_reduce_sa138 & multm_reduce_sd138;
  assign multm_reduce_add3b0_maj3b_wy139 = multm_reduce_sa139 & multm_reduce_sd139;
  assign multm_reduce_add3b0_maj3b_wy140 = multm_reduce_sa140 & multm_reduce_sd140;
  assign multm_reduce_add3b0_maj3b_wy141 = multm_reduce_sa141 & multm_reduce_sd141;
  assign multm_reduce_add3b0_maj3b_wy142 = multm_reduce_sa142 & multm_reduce_sd142;
  assign multm_reduce_add3b0_maj3b_wy143 = multm_reduce_sa143 & multm_reduce_sd143;
  assign multm_reduce_add3b0_maj3b_wy144 = multm_reduce_sa144 & multm_reduce_sd144;
  assign multm_reduce_add3b0_maj3b_wy145 = multm_reduce_sa145 & multm_reduce_sd145;
  assign multm_reduce_add3b0_maj3b_wy146 = multm_reduce_sa146 & multm_reduce_sd146;
  assign multm_reduce_add3b0_maj3b_wy147 = multm_reduce_sa147 & multm_reduce_sd147;
  assign multm_reduce_add3b0_maj3b_wy148 = multm_reduce_sa148 & multm_reduce_sd148;
  assign multm_reduce_add3b0_maj3b_wy149 = multm_reduce_sa149 & multm_reduce_sd149;
  assign multm_reduce_add3b0_maj3b_wy150 = multm_reduce_sa150 & multm_reduce_sd150;
  assign multm_reduce_add3b0_maj3b_wy151 = multm_reduce_sa151 & multm_reduce_sd151;
  assign multm_reduce_add3b0_maj3b_wy152 = multm_reduce_sa152 & multm_reduce_sd152;
  assign multm_reduce_add3b0_maj3b_wy153 = multm_reduce_sa153 & multm_reduce_sd153;
  assign multm_reduce_add3b0_maj3b_wy154 = multm_reduce_sa154 & multm_reduce_sd154;
  assign multm_reduce_add3b0_maj3b_wy155 = multm_reduce_sa155 & multm_reduce_sd155;
  assign multm_reduce_add3b0_maj3b_wy156 = multm_reduce_sa156 & multm_reduce_sd156;
  assign multm_reduce_add3b0_maj3b_wy157 = multm_reduce_sa157 & multm_reduce_sd157;
  assign multm_reduce_add3b0_maj3b_wy158 = multm_reduce_sa158 & multm_reduce_sd158;
  assign multm_reduce_add3b0_maj3b_wy159 = multm_reduce_sa159 & multm_reduce_sd159;
  assign multm_reduce_add3b0_maj3b_wy160 = multm_reduce_sa160 & multm_reduce_sd160;
  assign multm_reduce_add3b0_maj3b_wy161 = multm_reduce_sa161 & multm_reduce_sd161;
  assign multm_reduce_add3b0_maj3b_wy162 = multm_reduce_sa162 & multm_reduce_sd162;
  assign multm_reduce_add3b0_maj3b_wy163 = multm_reduce_sa163 & multm_reduce_sd163;
  assign multm_reduce_add3b0_maj3b_wy164 = multm_reduce_sa164 & multm_reduce_sd164;
  assign multm_reduce_add3b0_maj3b_wy165 = multm_reduce_sa165 & multm_reduce_sd165;
  assign multm_reduce_add3b0_maj3b_wy166 = multm_reduce_sa166 & multm_reduce_sd166;
  assign multm_reduce_add3b0_maj3b_wy167 = multm_reduce_sa167 & multm_reduce_sd167;
  assign multm_reduce_add3b0_maj3b_wy168 = multm_reduce_sa168 & multm_reduce_sd168;
  assign multm_reduce_add3b0_maj3b_wy169 = multm_reduce_sa169 & multm_reduce_sd169;
  assign multm_reduce_add3b0_maj3b_wy170 = multm_reduce_sa170 & multm_reduce_sd170;
  assign multm_reduce_add3b0_maj3b_wy171 = multm_reduce_sa171 & multm_reduce_sd171;
  assign multm_reduce_add3b0_maj3b_wy172 = multm_reduce_sa172 & multm_reduce_sd172;
  assign multm_reduce_add3b0_maj3b_wy173 = multm_reduce_sa173 & multm_reduce_sd173;
  assign multm_reduce_add3b0_maj3b_wy174 = multm_reduce_sa174 & multm_reduce_sd174;
  assign multm_reduce_add3b0_maj3b_wy175 = multm_reduce_sa175 & multm_reduce_sd175;
  assign multm_reduce_add3b0_maj3b_wy176 = multm_reduce_sa176 & multm_reduce_sd176;
  assign multm_reduce_add3b0_maj3b_wy177 = multm_reduce_sa177 & multm_reduce_sd177;
  assign multm_reduce_add3b0_maj3b_wy178 = multm_reduce_sa178 & multm_reduce_sd178;
  assign multm_reduce_add3b0_maj3b_wy179 = multm_reduce_sa179 & multm_reduce_sd179;
  assign multm_reduce_add3b0_maj3b_wy180 = multm_reduce_sa180 & multm_reduce_sd180;
  assign multm_reduce_add3b0_maj3b_wy181 = multm_reduce_sa181 & multm_reduce_sd181;
  assign multm_reduce_add3b0_maj3b_wy182 = multm_reduce_sa182 & multm_reduce_sd182;
  assign multm_reduce_add3b0_maj3b_xy0 = multm_reduce_sc0 & multm_reduce_sd0;
  assign multm_reduce_add3b0_maj3b_xy1 = multm_reduce_sc1 & multm_reduce_sd1;
  assign multm_reduce_add3b0_maj3b_xy2 = multm_reduce_sc2 & multm_reduce_sd2;
  assign multm_reduce_add3b0_maj3b_xy3 = multm_reduce_sc3 & multm_reduce_sd3;
  assign multm_reduce_add3b0_maj3b_xy4 = multm_reduce_sc4 & multm_reduce_sd4;
  assign multm_reduce_add3b0_maj3b_xy5 = multm_reduce_sc5 & multm_reduce_sd5;
  assign multm_reduce_add3b0_maj3b_xy6 = multm_reduce_sc6 & multm_reduce_sd6;
  assign multm_reduce_add3b0_maj3b_xy7 = multm_reduce_sc7 & multm_reduce_sd7;
  assign multm_reduce_add3b0_maj3b_xy8 = multm_reduce_sc8 & multm_reduce_sd8;
  assign multm_reduce_add3b0_maj3b_xy9 = multm_reduce_sc9 & multm_reduce_sd9;
  assign multm_reduce_add3b0_maj3b_xy10 = multm_reduce_sc10 & multm_reduce_sd10;
  assign multm_reduce_add3b0_maj3b_xy11 = multm_reduce_sc11 & multm_reduce_sd11;
  assign multm_reduce_add3b0_maj3b_xy12 = multm_reduce_sc12 & multm_reduce_sd12;
  assign multm_reduce_add3b0_maj3b_xy13 = multm_reduce_sc13 & multm_reduce_sd13;
  assign multm_reduce_add3b0_maj3b_xy14 = multm_reduce_sc14 & multm_reduce_sd14;
  assign multm_reduce_add3b0_maj3b_xy15 = multm_reduce_sc15 & multm_reduce_sd15;
  assign multm_reduce_add3b0_maj3b_xy16 = multm_reduce_sc16 & multm_reduce_sd16;
  assign multm_reduce_add3b0_maj3b_xy17 = multm_reduce_sc17 & multm_reduce_sd17;
  assign multm_reduce_add3b0_maj3b_xy18 = multm_reduce_sc18 & multm_reduce_sd18;
  assign multm_reduce_add3b0_maj3b_xy19 = multm_reduce_sc19 & multm_reduce_sd19;
  assign multm_reduce_add3b0_maj3b_xy20 = multm_reduce_sc20 & multm_reduce_sd20;
  assign multm_reduce_add3b0_maj3b_xy21 = multm_reduce_sc21 & multm_reduce_sd21;
  assign multm_reduce_add3b0_maj3b_xy22 = multm_reduce_sc22 & multm_reduce_sd22;
  assign multm_reduce_add3b0_maj3b_xy23 = multm_reduce_sc23 & multm_reduce_sd23;
  assign multm_reduce_add3b0_maj3b_xy24 = multm_reduce_sc24 & multm_reduce_sd24;
  assign multm_reduce_add3b0_maj3b_xy25 = multm_reduce_sc25 & multm_reduce_sd25;
  assign multm_reduce_add3b0_maj3b_xy26 = multm_reduce_sc26 & multm_reduce_sd26;
  assign multm_reduce_add3b0_maj3b_xy27 = multm_reduce_sc27 & multm_reduce_sd27;
  assign multm_reduce_add3b0_maj3b_xy28 = multm_reduce_sc28 & multm_reduce_sd28;
  assign multm_reduce_add3b0_maj3b_xy29 = multm_reduce_sc29 & multm_reduce_sd29;
  assign multm_reduce_add3b0_maj3b_xy30 = multm_reduce_sc30 & multm_reduce_sd30;
  assign multm_reduce_add3b0_maj3b_xy31 = multm_reduce_sc31 & multm_reduce_sd31;
  assign multm_reduce_add3b0_maj3b_xy32 = multm_reduce_sc32 & multm_reduce_sd32;
  assign multm_reduce_add3b0_maj3b_xy33 = multm_reduce_sc33 & multm_reduce_sd33;
  assign multm_reduce_add3b0_maj3b_xy34 = multm_reduce_sc34 & multm_reduce_sd34;
  assign multm_reduce_add3b0_maj3b_xy35 = multm_reduce_sc35 & multm_reduce_sd35;
  assign multm_reduce_add3b0_maj3b_xy36 = multm_reduce_sc36 & multm_reduce_sd36;
  assign multm_reduce_add3b0_maj3b_xy37 = multm_reduce_sc37 & multm_reduce_sd37;
  assign multm_reduce_add3b0_maj3b_xy38 = multm_reduce_sc38 & multm_reduce_sd38;
  assign multm_reduce_add3b0_maj3b_xy39 = multm_reduce_sc39 & multm_reduce_sd39;
  assign multm_reduce_add3b0_maj3b_xy40 = multm_reduce_sc40 & multm_reduce_sd40;
  assign multm_reduce_add3b0_maj3b_xy41 = multm_reduce_sc41 & multm_reduce_sd41;
  assign multm_reduce_add3b0_maj3b_xy42 = multm_reduce_sc42 & multm_reduce_sd42;
  assign multm_reduce_add3b0_maj3b_xy43 = multm_reduce_sc43 & multm_reduce_sd43;
  assign multm_reduce_add3b0_maj3b_xy44 = multm_reduce_sc44 & multm_reduce_sd44;
  assign multm_reduce_add3b0_maj3b_xy45 = multm_reduce_sc45 & multm_reduce_sd45;
  assign multm_reduce_add3b0_maj3b_xy46 = multm_reduce_sc46 & multm_reduce_sd46;
  assign multm_reduce_add3b0_maj3b_xy47 = multm_reduce_sc47 & multm_reduce_sd47;
  assign multm_reduce_add3b0_maj3b_xy48 = multm_reduce_sc48 & multm_reduce_sd48;
  assign multm_reduce_add3b0_maj3b_xy49 = multm_reduce_sc49 & multm_reduce_sd49;
  assign multm_reduce_add3b0_maj3b_xy50 = multm_reduce_sc50 & multm_reduce_sd50;
  assign multm_reduce_add3b0_maj3b_xy51 = multm_reduce_sc51 & multm_reduce_sd51;
  assign multm_reduce_add3b0_maj3b_xy52 = multm_reduce_sc52 & multm_reduce_sd52;
  assign multm_reduce_add3b0_maj3b_xy53 = multm_reduce_sc53 & multm_reduce_sd53;
  assign multm_reduce_add3b0_maj3b_xy54 = multm_reduce_sc54 & multm_reduce_sd54;
  assign multm_reduce_add3b0_maj3b_xy55 = multm_reduce_sc55 & multm_reduce_sd55;
  assign multm_reduce_add3b0_maj3b_xy56 = multm_reduce_sc56 & multm_reduce_sd56;
  assign multm_reduce_add3b0_maj3b_xy57 = multm_reduce_sc57 & multm_reduce_sd57;
  assign multm_reduce_add3b0_maj3b_xy58 = multm_reduce_sc58 & multm_reduce_sd58;
  assign multm_reduce_add3b0_maj3b_xy59 = multm_reduce_sc59 & multm_reduce_sd59;
  assign multm_reduce_add3b0_maj3b_xy60 = multm_reduce_sc60 & multm_reduce_sd60;
  assign multm_reduce_add3b0_maj3b_xy61 = multm_reduce_sc61 & multm_reduce_sd61;
  assign multm_reduce_add3b0_maj3b_xy62 = multm_reduce_sc62 & multm_reduce_sd62;
  assign multm_reduce_add3b0_maj3b_xy63 = multm_reduce_sc63 & multm_reduce_sd63;
  assign multm_reduce_add3b0_maj3b_xy64 = multm_reduce_sc64 & multm_reduce_sd64;
  assign multm_reduce_add3b0_maj3b_xy65 = multm_reduce_sc65 & multm_reduce_sd65;
  assign multm_reduce_add3b0_maj3b_xy66 = multm_reduce_sc66 & multm_reduce_sd66;
  assign multm_reduce_add3b0_maj3b_xy67 = multm_reduce_sc67 & multm_reduce_sd67;
  assign multm_reduce_add3b0_maj3b_xy68 = multm_reduce_sc68 & multm_reduce_sd68;
  assign multm_reduce_add3b0_maj3b_xy69 = multm_reduce_sc69 & multm_reduce_sd69;
  assign multm_reduce_add3b0_maj3b_xy70 = multm_reduce_sc70 & multm_reduce_sd70;
  assign multm_reduce_add3b0_maj3b_xy71 = multm_reduce_sc71 & multm_reduce_sd71;
  assign multm_reduce_add3b0_maj3b_xy72 = multm_reduce_sc72 & multm_reduce_sd72;
  assign multm_reduce_add3b0_maj3b_xy73 = multm_reduce_sc73 & multm_reduce_sd73;
  assign multm_reduce_add3b0_maj3b_xy74 = multm_reduce_sc74 & multm_reduce_sd74;
  assign multm_reduce_add3b0_maj3b_xy75 = multm_reduce_sc75 & multm_reduce_sd75;
  assign multm_reduce_add3b0_maj3b_xy76 = multm_reduce_sc76 & multm_reduce_sd76;
  assign multm_reduce_add3b0_maj3b_xy77 = multm_reduce_sc77 & multm_reduce_sd77;
  assign multm_reduce_add3b0_maj3b_xy78 = multm_reduce_sc78 & multm_reduce_sd78;
  assign multm_reduce_add3b0_maj3b_xy79 = multm_reduce_sc79 & multm_reduce_sd79;
  assign multm_reduce_add3b0_maj3b_xy80 = multm_reduce_sc80 & multm_reduce_sd80;
  assign multm_reduce_add3b0_maj3b_xy81 = multm_reduce_sc81 & multm_reduce_sd81;
  assign multm_reduce_add3b0_maj3b_xy82 = multm_reduce_sc82 & multm_reduce_sd82;
  assign multm_reduce_add3b0_maj3b_xy83 = multm_reduce_sc83 & multm_reduce_sd83;
  assign multm_reduce_add3b0_maj3b_xy84 = multm_reduce_sc84 & multm_reduce_sd84;
  assign multm_reduce_add3b0_maj3b_xy85 = multm_reduce_sc85 & multm_reduce_sd85;
  assign multm_reduce_add3b0_maj3b_xy86 = multm_reduce_sc86 & multm_reduce_sd86;
  assign multm_reduce_add3b0_maj3b_xy87 = multm_reduce_sc87 & multm_reduce_sd87;
  assign multm_reduce_add3b0_maj3b_xy88 = multm_reduce_sc88 & multm_reduce_sd88;
  assign multm_reduce_add3b0_maj3b_xy89 = multm_reduce_sc89 & multm_reduce_sd89;
  assign multm_reduce_add3b0_maj3b_xy90 = multm_reduce_sc90 & multm_reduce_sd90;
  assign multm_reduce_add3b0_maj3b_xy91 = multm_reduce_sc91 & multm_reduce_sd91;
  assign multm_reduce_add3b0_maj3b_xy92 = multm_reduce_sc92 & multm_reduce_sd92;
  assign multm_reduce_add3b0_maj3b_xy93 = multm_reduce_sc93 & multm_reduce_sd93;
  assign multm_reduce_add3b0_maj3b_xy94 = multm_reduce_sc94 & multm_reduce_sd94;
  assign multm_reduce_add3b0_maj3b_xy95 = multm_reduce_sc95 & multm_reduce_sd95;
  assign multm_reduce_add3b0_maj3b_xy96 = multm_reduce_sc96 & multm_reduce_sd96;
  assign multm_reduce_add3b0_maj3b_xy97 = multm_reduce_sc97 & multm_reduce_sd97;
  assign multm_reduce_add3b0_maj3b_xy98 = multm_reduce_sc98 & multm_reduce_sd98;
  assign multm_reduce_add3b0_maj3b_xy99 = multm_reduce_sc99 & multm_reduce_sd99;
  assign multm_reduce_add3b0_maj3b_xy100 = multm_reduce_sc100 & multm_reduce_sd100;
  assign multm_reduce_add3b0_maj3b_xy101 = multm_reduce_sc101 & multm_reduce_sd101;
  assign multm_reduce_add3b0_maj3b_xy102 = multm_reduce_sc102 & multm_reduce_sd102;
  assign multm_reduce_add3b0_maj3b_xy103 = multm_reduce_sc103 & multm_reduce_sd103;
  assign multm_reduce_add3b0_maj3b_xy104 = multm_reduce_sc104 & multm_reduce_sd104;
  assign multm_reduce_add3b0_maj3b_xy105 = multm_reduce_sc105 & multm_reduce_sd105;
  assign multm_reduce_add3b0_maj3b_xy106 = multm_reduce_sc106 & multm_reduce_sd106;
  assign multm_reduce_add3b0_maj3b_xy107 = multm_reduce_sc107 & multm_reduce_sd107;
  assign multm_reduce_add3b0_maj3b_xy108 = multm_reduce_sc108 & multm_reduce_sd108;
  assign multm_reduce_add3b0_maj3b_xy109 = multm_reduce_sc109 & multm_reduce_sd109;
  assign multm_reduce_add3b0_maj3b_xy110 = multm_reduce_sc110 & multm_reduce_sd110;
  assign multm_reduce_add3b0_maj3b_xy111 = multm_reduce_sc111 & multm_reduce_sd111;
  assign multm_reduce_add3b0_maj3b_xy112 = multm_reduce_sc112 & multm_reduce_sd112;
  assign multm_reduce_add3b0_maj3b_xy113 = multm_reduce_sc113 & multm_reduce_sd113;
  assign multm_reduce_add3b0_maj3b_xy114 = multm_reduce_sc114 & multm_reduce_sd114;
  assign multm_reduce_add3b0_maj3b_xy115 = multm_reduce_sc115 & multm_reduce_sd115;
  assign multm_reduce_add3b0_maj3b_xy116 = multm_reduce_sc116 & multm_reduce_sd116;
  assign multm_reduce_add3b0_maj3b_xy117 = multm_reduce_sc117 & multm_reduce_sd117;
  assign multm_reduce_add3b0_maj3b_xy118 = multm_reduce_sc118 & multm_reduce_sd118;
  assign multm_reduce_add3b0_maj3b_xy119 = multm_reduce_sc119 & multm_reduce_sd119;
  assign multm_reduce_add3b0_maj3b_xy120 = multm_reduce_sc120 & multm_reduce_sd120;
  assign multm_reduce_add3b0_maj3b_xy121 = multm_reduce_sc121 & multm_reduce_sd121;
  assign multm_reduce_add3b0_maj3b_xy122 = multm_reduce_sc122 & multm_reduce_sd122;
  assign multm_reduce_add3b0_maj3b_xy123 = multm_reduce_sc123 & multm_reduce_sd123;
  assign multm_reduce_add3b0_maj3b_xy124 = multm_reduce_sc124 & multm_reduce_sd124;
  assign multm_reduce_add3b0_maj3b_xy125 = multm_reduce_sc125 & multm_reduce_sd125;
  assign multm_reduce_add3b0_maj3b_xy126 = multm_reduce_sc126 & multm_reduce_sd126;
  assign multm_reduce_add3b0_maj3b_xy127 = multm_reduce_sc127 & multm_reduce_sd127;
  assign multm_reduce_add3b0_maj3b_xy128 = multm_reduce_sc128 & multm_reduce_sd128;
  assign multm_reduce_add3b0_maj3b_xy129 = multm_reduce_sc129 & multm_reduce_sd129;
  assign multm_reduce_add3b0_maj3b_xy130 = multm_reduce_sc130 & multm_reduce_sd130;
  assign multm_reduce_add3b0_maj3b_xy131 = multm_reduce_sc131 & multm_reduce_sd131;
  assign multm_reduce_add3b0_maj3b_xy132 = multm_reduce_sc132 & multm_reduce_sd132;
  assign multm_reduce_add3b0_maj3b_xy133 = multm_reduce_sc133 & multm_reduce_sd133;
  assign multm_reduce_add3b0_maj3b_xy134 = multm_reduce_sc134 & multm_reduce_sd134;
  assign multm_reduce_add3b0_maj3b_xy135 = multm_reduce_sc135 & multm_reduce_sd135;
  assign multm_reduce_add3b0_maj3b_xy136 = multm_reduce_sc136 & multm_reduce_sd136;
  assign multm_reduce_add3b0_maj3b_xy137 = multm_reduce_sc137 & multm_reduce_sd137;
  assign multm_reduce_add3b0_maj3b_xy138 = multm_reduce_sc138 & multm_reduce_sd138;
  assign multm_reduce_add3b0_maj3b_xy139 = multm_reduce_sc139 & multm_reduce_sd139;
  assign multm_reduce_add3b0_maj3b_xy140 = multm_reduce_sc140 & multm_reduce_sd140;
  assign multm_reduce_add3b0_maj3b_xy141 = multm_reduce_sc141 & multm_reduce_sd141;
  assign multm_reduce_add3b0_maj3b_xy142 = multm_reduce_sc142 & multm_reduce_sd142;
  assign multm_reduce_add3b0_maj3b_xy143 = multm_reduce_sc143 & multm_reduce_sd143;
  assign multm_reduce_add3b0_maj3b_xy144 = multm_reduce_sc144 & multm_reduce_sd144;
  assign multm_reduce_add3b0_maj3b_xy145 = multm_reduce_sc145 & multm_reduce_sd145;
  assign multm_reduce_add3b0_maj3b_xy146 = multm_reduce_sc146 & multm_reduce_sd146;
  assign multm_reduce_add3b0_maj3b_xy147 = multm_reduce_sc147 & multm_reduce_sd147;
  assign multm_reduce_add3b0_maj3b_xy148 = multm_reduce_sc148 & multm_reduce_sd148;
  assign multm_reduce_add3b0_maj3b_xy149 = multm_reduce_sc149 & multm_reduce_sd149;
  assign multm_reduce_add3b0_maj3b_xy150 = multm_reduce_sc150 & multm_reduce_sd150;
  assign multm_reduce_add3b0_maj3b_xy151 = multm_reduce_sc151 & multm_reduce_sd151;
  assign multm_reduce_add3b0_maj3b_xy152 = multm_reduce_sc152 & multm_reduce_sd152;
  assign multm_reduce_add3b0_maj3b_xy153 = multm_reduce_sc153 & multm_reduce_sd153;
  assign multm_reduce_add3b0_maj3b_xy154 = multm_reduce_sc154 & multm_reduce_sd154;
  assign multm_reduce_add3b0_maj3b_xy155 = multm_reduce_sc155 & multm_reduce_sd155;
  assign multm_reduce_add3b0_maj3b_xy156 = multm_reduce_sc156 & multm_reduce_sd156;
  assign multm_reduce_add3b0_maj3b_xy157 = multm_reduce_sc157 & multm_reduce_sd157;
  assign multm_reduce_add3b0_maj3b_xy158 = multm_reduce_sc158 & multm_reduce_sd158;
  assign multm_reduce_add3b0_maj3b_xy159 = multm_reduce_sc159 & multm_reduce_sd159;
  assign multm_reduce_add3b0_maj3b_xy160 = multm_reduce_sc160 & multm_reduce_sd160;
  assign multm_reduce_add3b0_maj3b_xy161 = multm_reduce_sc161 & multm_reduce_sd161;
  assign multm_reduce_add3b0_maj3b_xy162 = multm_reduce_sc162 & multm_reduce_sd162;
  assign multm_reduce_add3b0_maj3b_xy163 = multm_reduce_sc163 & multm_reduce_sd163;
  assign multm_reduce_add3b0_maj3b_xy164 = multm_reduce_sc164 & multm_reduce_sd164;
  assign multm_reduce_add3b0_maj3b_xy165 = multm_reduce_sc165 & multm_reduce_sd165;
  assign multm_reduce_add3b0_maj3b_xy166 = multm_reduce_sc166 & multm_reduce_sd166;
  assign multm_reduce_add3b0_maj3b_xy167 = multm_reduce_sc167 & multm_reduce_sd167;
  assign multm_reduce_add3b0_maj3b_xy168 = multm_reduce_sc168 & multm_reduce_sd168;
  assign multm_reduce_add3b0_maj3b_xy169 = multm_reduce_sc169 & multm_reduce_sd169;
  assign multm_reduce_add3b0_maj3b_xy170 = multm_reduce_sc170 & multm_reduce_sd170;
  assign multm_reduce_add3b0_maj3b_xy171 = multm_reduce_sc171 & multm_reduce_sd171;
  assign multm_reduce_add3b0_maj3b_xy172 = multm_reduce_sc172 & multm_reduce_sd172;
  assign multm_reduce_add3b0_maj3b_xy173 = multm_reduce_sc173 & multm_reduce_sd173;
  assign multm_reduce_add3b0_maj3b_xy174 = multm_reduce_sc174 & multm_reduce_sd174;
  assign multm_reduce_add3b0_maj3b_xy175 = multm_reduce_sc175 & multm_reduce_sd175;
  assign multm_reduce_add3b0_maj3b_xy176 = multm_reduce_sc176 & multm_reduce_sd176;
  assign multm_reduce_add3b0_maj3b_xy177 = multm_reduce_sc177 & multm_reduce_sd177;
  assign multm_reduce_add3b0_maj3b_xy178 = multm_reduce_sc178 & multm_reduce_sd178;
  assign multm_reduce_add3b0_maj3b_xy179 = multm_reduce_sc179 & multm_reduce_sd179;
  assign multm_reduce_add3b0_maj3b_xy180 = multm_reduce_sc180 & multm_reduce_sd180;
  assign multm_reduce_add3b0_maj3b_xy181 = multm_reduce_sc181 & multm_reduce_sd181;
  assign multm_reduce_add3b0_maj3b_xy182 = multm_reduce_sc182 & multm_reduce_sd182;
  assign multm_reduce_add3b0_xor3b_wx0 = multm_reduce_sa0 ^ multm_reduce_sc0;
  assign multm_reduce_add3b0_xor3b_wx1 = multm_reduce_sa1 ^ multm_reduce_sc1;
  assign multm_reduce_add3b0_xor3b_wx2 = multm_reduce_sa2 ^ multm_reduce_sc2;
  assign multm_reduce_add3b0_xor3b_wx3 = multm_reduce_sa3 ^ multm_reduce_sc3;
  assign multm_reduce_add3b0_xor3b_wx4 = multm_reduce_sa4 ^ multm_reduce_sc4;
  assign multm_reduce_add3b0_xor3b_wx5 = multm_reduce_sa5 ^ multm_reduce_sc5;
  assign multm_reduce_add3b0_xor3b_wx6 = multm_reduce_sa6 ^ multm_reduce_sc6;
  assign multm_reduce_add3b0_xor3b_wx7 = multm_reduce_sa7 ^ multm_reduce_sc7;
  assign multm_reduce_add3b0_xor3b_wx8 = multm_reduce_sa8 ^ multm_reduce_sc8;
  assign multm_reduce_add3b0_xor3b_wx9 = multm_reduce_sa9 ^ multm_reduce_sc9;
  assign multm_reduce_add3b0_xor3b_wx10 = multm_reduce_sa10 ^ multm_reduce_sc10;
  assign multm_reduce_add3b0_xor3b_wx11 = multm_reduce_sa11 ^ multm_reduce_sc11;
  assign multm_reduce_add3b0_xor3b_wx12 = multm_reduce_sa12 ^ multm_reduce_sc12;
  assign multm_reduce_add3b0_xor3b_wx13 = multm_reduce_sa13 ^ multm_reduce_sc13;
  assign multm_reduce_add3b0_xor3b_wx14 = multm_reduce_sa14 ^ multm_reduce_sc14;
  assign multm_reduce_add3b0_xor3b_wx15 = multm_reduce_sa15 ^ multm_reduce_sc15;
  assign multm_reduce_add3b0_xor3b_wx16 = multm_reduce_sa16 ^ multm_reduce_sc16;
  assign multm_reduce_add3b0_xor3b_wx17 = multm_reduce_sa17 ^ multm_reduce_sc17;
  assign multm_reduce_add3b0_xor3b_wx18 = multm_reduce_sa18 ^ multm_reduce_sc18;
  assign multm_reduce_add3b0_xor3b_wx19 = multm_reduce_sa19 ^ multm_reduce_sc19;
  assign multm_reduce_add3b0_xor3b_wx20 = multm_reduce_sa20 ^ multm_reduce_sc20;
  assign multm_reduce_add3b0_xor3b_wx21 = multm_reduce_sa21 ^ multm_reduce_sc21;
  assign multm_reduce_add3b0_xor3b_wx22 = multm_reduce_sa22 ^ multm_reduce_sc22;
  assign multm_reduce_add3b0_xor3b_wx23 = multm_reduce_sa23 ^ multm_reduce_sc23;
  assign multm_reduce_add3b0_xor3b_wx24 = multm_reduce_sa24 ^ multm_reduce_sc24;
  assign multm_reduce_add3b0_xor3b_wx25 = multm_reduce_sa25 ^ multm_reduce_sc25;
  assign multm_reduce_add3b0_xor3b_wx26 = multm_reduce_sa26 ^ multm_reduce_sc26;
  assign multm_reduce_add3b0_xor3b_wx27 = multm_reduce_sa27 ^ multm_reduce_sc27;
  assign multm_reduce_add3b0_xor3b_wx28 = multm_reduce_sa28 ^ multm_reduce_sc28;
  assign multm_reduce_add3b0_xor3b_wx29 = multm_reduce_sa29 ^ multm_reduce_sc29;
  assign multm_reduce_add3b0_xor3b_wx30 = multm_reduce_sa30 ^ multm_reduce_sc30;
  assign multm_reduce_add3b0_xor3b_wx31 = multm_reduce_sa31 ^ multm_reduce_sc31;
  assign multm_reduce_add3b0_xor3b_wx32 = multm_reduce_sa32 ^ multm_reduce_sc32;
  assign multm_reduce_add3b0_xor3b_wx33 = multm_reduce_sa33 ^ multm_reduce_sc33;
  assign multm_reduce_add3b0_xor3b_wx34 = multm_reduce_sa34 ^ multm_reduce_sc34;
  assign multm_reduce_add3b0_xor3b_wx35 = multm_reduce_sa35 ^ multm_reduce_sc35;
  assign multm_reduce_add3b0_xor3b_wx36 = multm_reduce_sa36 ^ multm_reduce_sc36;
  assign multm_reduce_add3b0_xor3b_wx37 = multm_reduce_sa37 ^ multm_reduce_sc37;
  assign multm_reduce_add3b0_xor3b_wx38 = multm_reduce_sa38 ^ multm_reduce_sc38;
  assign multm_reduce_add3b0_xor3b_wx39 = multm_reduce_sa39 ^ multm_reduce_sc39;
  assign multm_reduce_add3b0_xor3b_wx40 = multm_reduce_sa40 ^ multm_reduce_sc40;
  assign multm_reduce_add3b0_xor3b_wx41 = multm_reduce_sa41 ^ multm_reduce_sc41;
  assign multm_reduce_add3b0_xor3b_wx42 = multm_reduce_sa42 ^ multm_reduce_sc42;
  assign multm_reduce_add3b0_xor3b_wx43 = multm_reduce_sa43 ^ multm_reduce_sc43;
  assign multm_reduce_add3b0_xor3b_wx44 = multm_reduce_sa44 ^ multm_reduce_sc44;
  assign multm_reduce_add3b0_xor3b_wx45 = multm_reduce_sa45 ^ multm_reduce_sc45;
  assign multm_reduce_add3b0_xor3b_wx46 = multm_reduce_sa46 ^ multm_reduce_sc46;
  assign multm_reduce_add3b0_xor3b_wx47 = multm_reduce_sa47 ^ multm_reduce_sc47;
  assign multm_reduce_add3b0_xor3b_wx48 = multm_reduce_sa48 ^ multm_reduce_sc48;
  assign multm_reduce_add3b0_xor3b_wx49 = multm_reduce_sa49 ^ multm_reduce_sc49;
  assign multm_reduce_add3b0_xor3b_wx50 = multm_reduce_sa50 ^ multm_reduce_sc50;
  assign multm_reduce_add3b0_xor3b_wx51 = multm_reduce_sa51 ^ multm_reduce_sc51;
  assign multm_reduce_add3b0_xor3b_wx52 = multm_reduce_sa52 ^ multm_reduce_sc52;
  assign multm_reduce_add3b0_xor3b_wx53 = multm_reduce_sa53 ^ multm_reduce_sc53;
  assign multm_reduce_add3b0_xor3b_wx54 = multm_reduce_sa54 ^ multm_reduce_sc54;
  assign multm_reduce_add3b0_xor3b_wx55 = multm_reduce_sa55 ^ multm_reduce_sc55;
  assign multm_reduce_add3b0_xor3b_wx56 = multm_reduce_sa56 ^ multm_reduce_sc56;
  assign multm_reduce_add3b0_xor3b_wx57 = multm_reduce_sa57 ^ multm_reduce_sc57;
  assign multm_reduce_add3b0_xor3b_wx58 = multm_reduce_sa58 ^ multm_reduce_sc58;
  assign multm_reduce_add3b0_xor3b_wx59 = multm_reduce_sa59 ^ multm_reduce_sc59;
  assign multm_reduce_add3b0_xor3b_wx60 = multm_reduce_sa60 ^ multm_reduce_sc60;
  assign multm_reduce_add3b0_xor3b_wx61 = multm_reduce_sa61 ^ multm_reduce_sc61;
  assign multm_reduce_add3b0_xor3b_wx62 = multm_reduce_sa62 ^ multm_reduce_sc62;
  assign multm_reduce_add3b0_xor3b_wx63 = multm_reduce_sa63 ^ multm_reduce_sc63;
  assign multm_reduce_add3b0_xor3b_wx64 = multm_reduce_sa64 ^ multm_reduce_sc64;
  assign multm_reduce_add3b0_xor3b_wx65 = multm_reduce_sa65 ^ multm_reduce_sc65;
  assign multm_reduce_add3b0_xor3b_wx66 = multm_reduce_sa66 ^ multm_reduce_sc66;
  assign multm_reduce_add3b0_xor3b_wx67 = multm_reduce_sa67 ^ multm_reduce_sc67;
  assign multm_reduce_add3b0_xor3b_wx68 = multm_reduce_sa68 ^ multm_reduce_sc68;
  assign multm_reduce_add3b0_xor3b_wx69 = multm_reduce_sa69 ^ multm_reduce_sc69;
  assign multm_reduce_add3b0_xor3b_wx70 = multm_reduce_sa70 ^ multm_reduce_sc70;
  assign multm_reduce_add3b0_xor3b_wx71 = multm_reduce_sa71 ^ multm_reduce_sc71;
  assign multm_reduce_add3b0_xor3b_wx72 = multm_reduce_sa72 ^ multm_reduce_sc72;
  assign multm_reduce_add3b0_xor3b_wx73 = multm_reduce_sa73 ^ multm_reduce_sc73;
  assign multm_reduce_add3b0_xor3b_wx74 = multm_reduce_sa74 ^ multm_reduce_sc74;
  assign multm_reduce_add3b0_xor3b_wx75 = multm_reduce_sa75 ^ multm_reduce_sc75;
  assign multm_reduce_add3b0_xor3b_wx76 = multm_reduce_sa76 ^ multm_reduce_sc76;
  assign multm_reduce_add3b0_xor3b_wx77 = multm_reduce_sa77 ^ multm_reduce_sc77;
  assign multm_reduce_add3b0_xor3b_wx78 = multm_reduce_sa78 ^ multm_reduce_sc78;
  assign multm_reduce_add3b0_xor3b_wx79 = multm_reduce_sa79 ^ multm_reduce_sc79;
  assign multm_reduce_add3b0_xor3b_wx80 = multm_reduce_sa80 ^ multm_reduce_sc80;
  assign multm_reduce_add3b0_xor3b_wx81 = multm_reduce_sa81 ^ multm_reduce_sc81;
  assign multm_reduce_add3b0_xor3b_wx82 = multm_reduce_sa82 ^ multm_reduce_sc82;
  assign multm_reduce_add3b0_xor3b_wx83 = multm_reduce_sa83 ^ multm_reduce_sc83;
  assign multm_reduce_add3b0_xor3b_wx84 = multm_reduce_sa84 ^ multm_reduce_sc84;
  assign multm_reduce_add3b0_xor3b_wx85 = multm_reduce_sa85 ^ multm_reduce_sc85;
  assign multm_reduce_add3b0_xor3b_wx86 = multm_reduce_sa86 ^ multm_reduce_sc86;
  assign multm_reduce_add3b0_xor3b_wx87 = multm_reduce_sa87 ^ multm_reduce_sc87;
  assign multm_reduce_add3b0_xor3b_wx88 = multm_reduce_sa88 ^ multm_reduce_sc88;
  assign multm_reduce_add3b0_xor3b_wx89 = multm_reduce_sa89 ^ multm_reduce_sc89;
  assign multm_reduce_add3b0_xor3b_wx90 = multm_reduce_sa90 ^ multm_reduce_sc90;
  assign multm_reduce_add3b0_xor3b_wx91 = multm_reduce_sa91 ^ multm_reduce_sc91;
  assign multm_reduce_add3b0_xor3b_wx92 = multm_reduce_sa92 ^ multm_reduce_sc92;
  assign multm_reduce_add3b0_xor3b_wx93 = multm_reduce_sa93 ^ multm_reduce_sc93;
  assign multm_reduce_add3b0_xor3b_wx94 = multm_reduce_sa94 ^ multm_reduce_sc94;
  assign multm_reduce_add3b0_xor3b_wx95 = multm_reduce_sa95 ^ multm_reduce_sc95;
  assign multm_reduce_add3b0_xor3b_wx96 = multm_reduce_sa96 ^ multm_reduce_sc96;
  assign multm_reduce_add3b0_xor3b_wx97 = multm_reduce_sa97 ^ multm_reduce_sc97;
  assign multm_reduce_add3b0_xor3b_wx98 = multm_reduce_sa98 ^ multm_reduce_sc98;
  assign multm_reduce_add3b0_xor3b_wx99 = multm_reduce_sa99 ^ multm_reduce_sc99;
  assign multm_reduce_add3b0_xor3b_wx100 = multm_reduce_sa100 ^ multm_reduce_sc100;
  assign multm_reduce_add3b0_xor3b_wx101 = multm_reduce_sa101 ^ multm_reduce_sc101;
  assign multm_reduce_add3b0_xor3b_wx102 = multm_reduce_sa102 ^ multm_reduce_sc102;
  assign multm_reduce_add3b0_xor3b_wx103 = multm_reduce_sa103 ^ multm_reduce_sc103;
  assign multm_reduce_add3b0_xor3b_wx104 = multm_reduce_sa104 ^ multm_reduce_sc104;
  assign multm_reduce_add3b0_xor3b_wx105 = multm_reduce_sa105 ^ multm_reduce_sc105;
  assign multm_reduce_add3b0_xor3b_wx106 = multm_reduce_sa106 ^ multm_reduce_sc106;
  assign multm_reduce_add3b0_xor3b_wx107 = multm_reduce_sa107 ^ multm_reduce_sc107;
  assign multm_reduce_add3b0_xor3b_wx108 = multm_reduce_sa108 ^ multm_reduce_sc108;
  assign multm_reduce_add3b0_xor3b_wx109 = multm_reduce_sa109 ^ multm_reduce_sc109;
  assign multm_reduce_add3b0_xor3b_wx110 = multm_reduce_sa110 ^ multm_reduce_sc110;
  assign multm_reduce_add3b0_xor3b_wx111 = multm_reduce_sa111 ^ multm_reduce_sc111;
  assign multm_reduce_add3b0_xor3b_wx112 = multm_reduce_sa112 ^ multm_reduce_sc112;
  assign multm_reduce_add3b0_xor3b_wx113 = multm_reduce_sa113 ^ multm_reduce_sc113;
  assign multm_reduce_add3b0_xor3b_wx114 = multm_reduce_sa114 ^ multm_reduce_sc114;
  assign multm_reduce_add3b0_xor3b_wx115 = multm_reduce_sa115 ^ multm_reduce_sc115;
  assign multm_reduce_add3b0_xor3b_wx116 = multm_reduce_sa116 ^ multm_reduce_sc116;
  assign multm_reduce_add3b0_xor3b_wx117 = multm_reduce_sa117 ^ multm_reduce_sc117;
  assign multm_reduce_add3b0_xor3b_wx118 = multm_reduce_sa118 ^ multm_reduce_sc118;
  assign multm_reduce_add3b0_xor3b_wx119 = multm_reduce_sa119 ^ multm_reduce_sc119;
  assign multm_reduce_add3b0_xor3b_wx120 = multm_reduce_sa120 ^ multm_reduce_sc120;
  assign multm_reduce_add3b0_xor3b_wx121 = multm_reduce_sa121 ^ multm_reduce_sc121;
  assign multm_reduce_add3b0_xor3b_wx122 = multm_reduce_sa122 ^ multm_reduce_sc122;
  assign multm_reduce_add3b0_xor3b_wx123 = multm_reduce_sa123 ^ multm_reduce_sc123;
  assign multm_reduce_add3b0_xor3b_wx124 = multm_reduce_sa124 ^ multm_reduce_sc124;
  assign multm_reduce_add3b0_xor3b_wx125 = multm_reduce_sa125 ^ multm_reduce_sc125;
  assign multm_reduce_add3b0_xor3b_wx126 = multm_reduce_sa126 ^ multm_reduce_sc126;
  assign multm_reduce_add3b0_xor3b_wx127 = multm_reduce_sa127 ^ multm_reduce_sc127;
  assign multm_reduce_add3b0_xor3b_wx128 = multm_reduce_sa128 ^ multm_reduce_sc128;
  assign multm_reduce_add3b0_xor3b_wx129 = multm_reduce_sa129 ^ multm_reduce_sc129;
  assign multm_reduce_add3b0_xor3b_wx130 = multm_reduce_sa130 ^ multm_reduce_sc130;
  assign multm_reduce_add3b0_xor3b_wx131 = multm_reduce_sa131 ^ multm_reduce_sc131;
  assign multm_reduce_add3b0_xor3b_wx132 = multm_reduce_sa132 ^ multm_reduce_sc132;
  assign multm_reduce_add3b0_xor3b_wx133 = multm_reduce_sa133 ^ multm_reduce_sc133;
  assign multm_reduce_add3b0_xor3b_wx134 = multm_reduce_sa134 ^ multm_reduce_sc134;
  assign multm_reduce_add3b0_xor3b_wx135 = multm_reduce_sa135 ^ multm_reduce_sc135;
  assign multm_reduce_add3b0_xor3b_wx136 = multm_reduce_sa136 ^ multm_reduce_sc136;
  assign multm_reduce_add3b0_xor3b_wx137 = multm_reduce_sa137 ^ multm_reduce_sc137;
  assign multm_reduce_add3b0_xor3b_wx138 = multm_reduce_sa138 ^ multm_reduce_sc138;
  assign multm_reduce_add3b0_xor3b_wx139 = multm_reduce_sa139 ^ multm_reduce_sc139;
  assign multm_reduce_add3b0_xor3b_wx140 = multm_reduce_sa140 ^ multm_reduce_sc140;
  assign multm_reduce_add3b0_xor3b_wx141 = multm_reduce_sa141 ^ multm_reduce_sc141;
  assign multm_reduce_add3b0_xor3b_wx142 = multm_reduce_sa142 ^ multm_reduce_sc142;
  assign multm_reduce_add3b0_xor3b_wx143 = multm_reduce_sa143 ^ multm_reduce_sc143;
  assign multm_reduce_add3b0_xor3b_wx144 = multm_reduce_sa144 ^ multm_reduce_sc144;
  assign multm_reduce_add3b0_xor3b_wx145 = multm_reduce_sa145 ^ multm_reduce_sc145;
  assign multm_reduce_add3b0_xor3b_wx146 = multm_reduce_sa146 ^ multm_reduce_sc146;
  assign multm_reduce_add3b0_xor3b_wx147 = multm_reduce_sa147 ^ multm_reduce_sc147;
  assign multm_reduce_add3b0_xor3b_wx148 = multm_reduce_sa148 ^ multm_reduce_sc148;
  assign multm_reduce_add3b0_xor3b_wx149 = multm_reduce_sa149 ^ multm_reduce_sc149;
  assign multm_reduce_add3b0_xor3b_wx150 = multm_reduce_sa150 ^ multm_reduce_sc150;
  assign multm_reduce_add3b0_xor3b_wx151 = multm_reduce_sa151 ^ multm_reduce_sc151;
  assign multm_reduce_add3b0_xor3b_wx152 = multm_reduce_sa152 ^ multm_reduce_sc152;
  assign multm_reduce_add3b0_xor3b_wx153 = multm_reduce_sa153 ^ multm_reduce_sc153;
  assign multm_reduce_add3b0_xor3b_wx154 = multm_reduce_sa154 ^ multm_reduce_sc154;
  assign multm_reduce_add3b0_xor3b_wx155 = multm_reduce_sa155 ^ multm_reduce_sc155;
  assign multm_reduce_add3b0_xor3b_wx156 = multm_reduce_sa156 ^ multm_reduce_sc156;
  assign multm_reduce_add3b0_xor3b_wx157 = multm_reduce_sa157 ^ multm_reduce_sc157;
  assign multm_reduce_add3b0_xor3b_wx158 = multm_reduce_sa158 ^ multm_reduce_sc158;
  assign multm_reduce_add3b0_xor3b_wx159 = multm_reduce_sa159 ^ multm_reduce_sc159;
  assign multm_reduce_add3b0_xor3b_wx160 = multm_reduce_sa160 ^ multm_reduce_sc160;
  assign multm_reduce_add3b0_xor3b_wx161 = multm_reduce_sa161 ^ multm_reduce_sc161;
  assign multm_reduce_add3b0_xor3b_wx162 = multm_reduce_sa162 ^ multm_reduce_sc162;
  assign multm_reduce_add3b0_xor3b_wx163 = multm_reduce_sa163 ^ multm_reduce_sc163;
  assign multm_reduce_add3b0_xor3b_wx164 = multm_reduce_sa164 ^ multm_reduce_sc164;
  assign multm_reduce_add3b0_xor3b_wx165 = multm_reduce_sa165 ^ multm_reduce_sc165;
  assign multm_reduce_add3b0_xor3b_wx166 = multm_reduce_sa166 ^ multm_reduce_sc166;
  assign multm_reduce_add3b0_xor3b_wx167 = multm_reduce_sa167 ^ multm_reduce_sc167;
  assign multm_reduce_add3b0_xor3b_wx168 = multm_reduce_sa168 ^ multm_reduce_sc168;
  assign multm_reduce_add3b0_xor3b_wx169 = multm_reduce_sa169 ^ multm_reduce_sc169;
  assign multm_reduce_add3b0_xor3b_wx170 = multm_reduce_sa170 ^ multm_reduce_sc170;
  assign multm_reduce_add3b0_xor3b_wx171 = multm_reduce_sa171 ^ multm_reduce_sc171;
  assign multm_reduce_add3b0_xor3b_wx172 = multm_reduce_sa172 ^ multm_reduce_sc172;
  assign multm_reduce_add3b0_xor3b_wx173 = multm_reduce_sa173 ^ multm_reduce_sc173;
  assign multm_reduce_add3b0_xor3b_wx174 = multm_reduce_sa174 ^ multm_reduce_sc174;
  assign multm_reduce_add3b0_xor3b_wx175 = multm_reduce_sa175 ^ multm_reduce_sc175;
  assign multm_reduce_add3b0_xor3b_wx176 = multm_reduce_sa176 ^ multm_reduce_sc176;
  assign multm_reduce_add3b0_xor3b_wx177 = multm_reduce_sa177 ^ multm_reduce_sc177;
  assign multm_reduce_add3b0_xor3b_wx178 = multm_reduce_sa178 ^ multm_reduce_sc178;
  assign multm_reduce_add3b0_xor3b_wx179 = multm_reduce_sa179 ^ multm_reduce_sc179;
  assign multm_reduce_add3b0_xor3b_wx180 = multm_reduce_sa180 ^ multm_reduce_sc180;
  assign multm_reduce_add3b0_xor3b_wx181 = multm_reduce_sa181 ^ multm_reduce_sc181;
  assign multm_reduce_add3b0_xor3b_wx182 = multm_reduce_sa182 ^ multm_reduce_sc182;
  assign multm_reduce_add3b1_maj3b_or3b_wx0 = multm_reduce_add3b1_maj3b_wx0 | multm_reduce_add3b1_maj3b_wy0;
  assign multm_reduce_add3b1_maj3b_or3b_wx1 = multm_reduce_add3b1_maj3b_wx1 | multm_reduce_add3b1_maj3b_wy1;
  assign multm_reduce_add3b1_maj3b_or3b_wx2 = multm_reduce_add3b1_maj3b_wx2 | multm_reduce_add3b1_maj3b_wy2;
  assign multm_reduce_add3b1_maj3b_or3b_wx3 = multm_reduce_add3b1_maj3b_wx3 | multm_reduce_add3b1_maj3b_wy3;
  assign multm_reduce_add3b1_maj3b_or3b_wx4 = multm_reduce_add3b1_maj3b_wx4 | multm_reduce_add3b1_maj3b_wy4;
  assign multm_reduce_add3b1_maj3b_or3b_wx5 = multm_reduce_add3b1_maj3b_wx5 | multm_reduce_add3b1_maj3b_wy5;
  assign multm_reduce_add3b1_maj3b_or3b_wx6 = multm_reduce_add3b1_maj3b_wx6 | multm_reduce_add3b1_maj3b_wy6;
  assign multm_reduce_add3b1_maj3b_or3b_wx7 = multm_reduce_add3b1_maj3b_wx7 | multm_reduce_add3b1_maj3b_wy7;
  assign multm_reduce_add3b1_maj3b_or3b_wx8 = multm_reduce_add3b1_maj3b_wx8 | multm_reduce_add3b1_maj3b_wy8;
  assign multm_reduce_add3b1_maj3b_or3b_wx9 = multm_reduce_add3b1_maj3b_wx9 | multm_reduce_add3b1_maj3b_wy9;
  assign multm_reduce_add3b1_maj3b_or3b_wx10 = multm_reduce_add3b1_maj3b_wx10 | multm_reduce_add3b1_maj3b_wy10;
  assign multm_reduce_add3b1_maj3b_or3b_wx11 = multm_reduce_add3b1_maj3b_wx11 | multm_reduce_add3b1_maj3b_wy11;
  assign multm_reduce_add3b1_maj3b_or3b_wx12 = multm_reduce_add3b1_maj3b_wx12 | multm_reduce_add3b1_maj3b_wy12;
  assign multm_reduce_add3b1_maj3b_or3b_wx13 = multm_reduce_add3b1_maj3b_wx13 | multm_reduce_add3b1_maj3b_wy13;
  assign multm_reduce_add3b1_maj3b_or3b_wx14 = multm_reduce_add3b1_maj3b_wx14 | multm_reduce_add3b1_maj3b_wy14;
  assign multm_reduce_add3b1_maj3b_or3b_wx15 = multm_reduce_add3b1_maj3b_wx15 | multm_reduce_add3b1_maj3b_wy15;
  assign multm_reduce_add3b1_maj3b_or3b_wx16 = multm_reduce_add3b1_maj3b_wx16 | multm_reduce_add3b1_maj3b_wy16;
  assign multm_reduce_add3b1_maj3b_or3b_wx17 = multm_reduce_add3b1_maj3b_wx17 | multm_reduce_add3b1_maj3b_wy17;
  assign multm_reduce_add3b1_maj3b_or3b_wx18 = multm_reduce_add3b1_maj3b_wx18 | multm_reduce_add3b1_maj3b_wy18;
  assign multm_reduce_add3b1_maj3b_or3b_wx19 = multm_reduce_add3b1_maj3b_wx19 | multm_reduce_add3b1_maj3b_wy19;
  assign multm_reduce_add3b1_maj3b_or3b_wx20 = multm_reduce_add3b1_maj3b_wx20 | multm_reduce_add3b1_maj3b_wy20;
  assign multm_reduce_add3b1_maj3b_or3b_wx21 = multm_reduce_add3b1_maj3b_wx21 | multm_reduce_add3b1_maj3b_wy21;
  assign multm_reduce_add3b1_maj3b_or3b_wx22 = multm_reduce_add3b1_maj3b_wx22 | multm_reduce_add3b1_maj3b_wy22;
  assign multm_reduce_add3b1_maj3b_or3b_wx23 = multm_reduce_add3b1_maj3b_wx23 | multm_reduce_add3b1_maj3b_wy23;
  assign multm_reduce_add3b1_maj3b_or3b_wx24 = multm_reduce_add3b1_maj3b_wx24 | multm_reduce_add3b1_maj3b_wy24;
  assign multm_reduce_add3b1_maj3b_or3b_wx25 = multm_reduce_add3b1_maj3b_wx25 | multm_reduce_add3b1_maj3b_wy25;
  assign multm_reduce_add3b1_maj3b_or3b_wx26 = multm_reduce_add3b1_maj3b_wx26 | multm_reduce_add3b1_maj3b_wy26;
  assign multm_reduce_add3b1_maj3b_or3b_wx27 = multm_reduce_add3b1_maj3b_wx27 | multm_reduce_add3b1_maj3b_wy27;
  assign multm_reduce_add3b1_maj3b_or3b_wx28 = multm_reduce_add3b1_maj3b_wx28 | multm_reduce_add3b1_maj3b_wy28;
  assign multm_reduce_add3b1_maj3b_or3b_wx29 = multm_reduce_add3b1_maj3b_wx29 | multm_reduce_add3b1_maj3b_wy29;
  assign multm_reduce_add3b1_maj3b_or3b_wx30 = multm_reduce_add3b1_maj3b_wx30 | multm_reduce_add3b1_maj3b_wy30;
  assign multm_reduce_add3b1_maj3b_or3b_wx31 = multm_reduce_add3b1_maj3b_wx31 | multm_reduce_add3b1_maj3b_wy31;
  assign multm_reduce_add3b1_maj3b_or3b_wx32 = multm_reduce_add3b1_maj3b_wx32 | multm_reduce_add3b1_maj3b_wy32;
  assign multm_reduce_add3b1_maj3b_or3b_wx33 = multm_reduce_add3b1_maj3b_wx33 | multm_reduce_add3b1_maj3b_wy33;
  assign multm_reduce_add3b1_maj3b_or3b_wx34 = multm_reduce_add3b1_maj3b_wx34 | multm_reduce_add3b1_maj3b_wy34;
  assign multm_reduce_add3b1_maj3b_or3b_wx35 = multm_reduce_add3b1_maj3b_wx35 | multm_reduce_add3b1_maj3b_wy35;
  assign multm_reduce_add3b1_maj3b_or3b_wx36 = multm_reduce_add3b1_maj3b_wx36 | multm_reduce_add3b1_maj3b_wy36;
  assign multm_reduce_add3b1_maj3b_or3b_wx37 = multm_reduce_add3b1_maj3b_wx37 | multm_reduce_add3b1_maj3b_wy37;
  assign multm_reduce_add3b1_maj3b_or3b_wx38 = multm_reduce_add3b1_maj3b_wx38 | multm_reduce_add3b1_maj3b_wy38;
  assign multm_reduce_add3b1_maj3b_or3b_wx39 = multm_reduce_add3b1_maj3b_wx39 | multm_reduce_add3b1_maj3b_wy39;
  assign multm_reduce_add3b1_maj3b_or3b_wx40 = multm_reduce_add3b1_maj3b_wx40 | multm_reduce_add3b1_maj3b_wy40;
  assign multm_reduce_add3b1_maj3b_or3b_wx41 = multm_reduce_add3b1_maj3b_wx41 | multm_reduce_add3b1_maj3b_wy41;
  assign multm_reduce_add3b1_maj3b_or3b_wx42 = multm_reduce_add3b1_maj3b_wx42 | multm_reduce_add3b1_maj3b_wy42;
  assign multm_reduce_add3b1_maj3b_or3b_wx43 = multm_reduce_add3b1_maj3b_wx43 | multm_reduce_add3b1_maj3b_wy43;
  assign multm_reduce_add3b1_maj3b_or3b_wx44 = multm_reduce_add3b1_maj3b_wx44 | multm_reduce_add3b1_maj3b_wy44;
  assign multm_reduce_add3b1_maj3b_or3b_wx45 = multm_reduce_add3b1_maj3b_wx45 | multm_reduce_add3b1_maj3b_wy45;
  assign multm_reduce_add3b1_maj3b_or3b_wx46 = multm_reduce_add3b1_maj3b_wx46 | multm_reduce_add3b1_maj3b_wy46;
  assign multm_reduce_add3b1_maj3b_or3b_wx47 = multm_reduce_add3b1_maj3b_wx47 | multm_reduce_add3b1_maj3b_wy47;
  assign multm_reduce_add3b1_maj3b_or3b_wx48 = multm_reduce_add3b1_maj3b_wx48 | multm_reduce_add3b1_maj3b_wy48;
  assign multm_reduce_add3b1_maj3b_or3b_wx49 = multm_reduce_add3b1_maj3b_wx49 | multm_reduce_add3b1_maj3b_wy49;
  assign multm_reduce_add3b1_maj3b_or3b_wx50 = multm_reduce_add3b1_maj3b_wx50 | multm_reduce_add3b1_maj3b_wy50;
  assign multm_reduce_add3b1_maj3b_or3b_wx51 = multm_reduce_add3b1_maj3b_wx51 | multm_reduce_add3b1_maj3b_wy51;
  assign multm_reduce_add3b1_maj3b_or3b_wx52 = multm_reduce_add3b1_maj3b_wx52 | multm_reduce_add3b1_maj3b_wy52;
  assign multm_reduce_add3b1_maj3b_or3b_wx53 = multm_reduce_add3b1_maj3b_wx53 | multm_reduce_add3b1_maj3b_wy53;
  assign multm_reduce_add3b1_maj3b_or3b_wx54 = multm_reduce_add3b1_maj3b_wx54 | multm_reduce_add3b1_maj3b_wy54;
  assign multm_reduce_add3b1_maj3b_or3b_wx55 = multm_reduce_add3b1_maj3b_wx55 | multm_reduce_add3b1_maj3b_wy55;
  assign multm_reduce_add3b1_maj3b_or3b_wx56 = multm_reduce_add3b1_maj3b_wx56 | multm_reduce_add3b1_maj3b_wy56;
  assign multm_reduce_add3b1_maj3b_or3b_wx57 = multm_reduce_add3b1_maj3b_wx57 | multm_reduce_add3b1_maj3b_wy57;
  assign multm_reduce_add3b1_maj3b_or3b_wx58 = multm_reduce_add3b1_maj3b_wx58 | multm_reduce_add3b1_maj3b_wy58;
  assign multm_reduce_add3b1_maj3b_or3b_wx59 = multm_reduce_add3b1_maj3b_wx59 | multm_reduce_add3b1_maj3b_wy59;
  assign multm_reduce_add3b1_maj3b_or3b_wx60 = multm_reduce_add3b1_maj3b_wx60 | multm_reduce_add3b1_maj3b_wy60;
  assign multm_reduce_add3b1_maj3b_or3b_wx61 = multm_reduce_add3b1_maj3b_wx61 | multm_reduce_add3b1_maj3b_wy61;
  assign multm_reduce_add3b1_maj3b_or3b_wx62 = multm_reduce_add3b1_maj3b_wx62 | multm_reduce_add3b1_maj3b_wy62;
  assign multm_reduce_add3b1_maj3b_or3b_wx63 = multm_reduce_add3b1_maj3b_wx63 | multm_reduce_add3b1_maj3b_wy63;
  assign multm_reduce_add3b1_maj3b_or3b_wx64 = multm_reduce_add3b1_maj3b_wx64 | multm_reduce_add3b1_maj3b_wy64;
  assign multm_reduce_add3b1_maj3b_or3b_wx65 = multm_reduce_add3b1_maj3b_wx65 | multm_reduce_add3b1_maj3b_wy65;
  assign multm_reduce_add3b1_maj3b_or3b_wx66 = multm_reduce_add3b1_maj3b_wx66 | multm_reduce_add3b1_maj3b_wy66;
  assign multm_reduce_add3b1_maj3b_or3b_wx67 = multm_reduce_add3b1_maj3b_wx67 | multm_reduce_add3b1_maj3b_wy67;
  assign multm_reduce_add3b1_maj3b_or3b_wx68 = multm_reduce_add3b1_maj3b_wx68 | multm_reduce_add3b1_maj3b_wy68;
  assign multm_reduce_add3b1_maj3b_or3b_wx69 = multm_reduce_add3b1_maj3b_wx69 | multm_reduce_add3b1_maj3b_wy69;
  assign multm_reduce_add3b1_maj3b_or3b_wx70 = multm_reduce_add3b1_maj3b_wx70 | multm_reduce_add3b1_maj3b_wy70;
  assign multm_reduce_add3b1_maj3b_or3b_wx71 = multm_reduce_add3b1_maj3b_wx71 | multm_reduce_add3b1_maj3b_wy71;
  assign multm_reduce_add3b1_maj3b_or3b_wx72 = multm_reduce_add3b1_maj3b_wx72 | multm_reduce_add3b1_maj3b_wy72;
  assign multm_reduce_add3b1_maj3b_or3b_wx73 = multm_reduce_add3b1_maj3b_wx73 | multm_reduce_add3b1_maj3b_wy73;
  assign multm_reduce_add3b1_maj3b_or3b_wx74 = multm_reduce_add3b1_maj3b_wx74 | multm_reduce_add3b1_maj3b_wy74;
  assign multm_reduce_add3b1_maj3b_or3b_wx75 = multm_reduce_add3b1_maj3b_wx75 | multm_reduce_add3b1_maj3b_wy75;
  assign multm_reduce_add3b1_maj3b_or3b_wx76 = multm_reduce_add3b1_maj3b_wx76 | multm_reduce_add3b1_maj3b_wy76;
  assign multm_reduce_add3b1_maj3b_or3b_wx77 = multm_reduce_add3b1_maj3b_wx77 | multm_reduce_add3b1_maj3b_wy77;
  assign multm_reduce_add3b1_maj3b_or3b_wx78 = multm_reduce_add3b1_maj3b_wx78 | multm_reduce_add3b1_maj3b_wy78;
  assign multm_reduce_add3b1_maj3b_or3b_wx79 = multm_reduce_add3b1_maj3b_wx79 | multm_reduce_add3b1_maj3b_wy79;
  assign multm_reduce_add3b1_maj3b_or3b_wx80 = multm_reduce_add3b1_maj3b_wx80 | multm_reduce_add3b1_maj3b_wy80;
  assign multm_reduce_add3b1_maj3b_or3b_wx81 = multm_reduce_add3b1_maj3b_wx81 | multm_reduce_add3b1_maj3b_wy81;
  assign multm_reduce_add3b1_maj3b_or3b_wx82 = multm_reduce_add3b1_maj3b_wx82 | multm_reduce_add3b1_maj3b_wy82;
  assign multm_reduce_add3b1_maj3b_or3b_wx83 = multm_reduce_add3b1_maj3b_wx83 | multm_reduce_add3b1_maj3b_wy83;
  assign multm_reduce_add3b1_maj3b_or3b_wx84 = multm_reduce_add3b1_maj3b_wx84 | multm_reduce_add3b1_maj3b_wy84;
  assign multm_reduce_add3b1_maj3b_or3b_wx85 = multm_reduce_add3b1_maj3b_wx85 | multm_reduce_add3b1_maj3b_wy85;
  assign multm_reduce_add3b1_maj3b_or3b_wx86 = multm_reduce_add3b1_maj3b_wx86 | multm_reduce_add3b1_maj3b_wy86;
  assign multm_reduce_add3b1_maj3b_or3b_wx87 = multm_reduce_add3b1_maj3b_wx87 | multm_reduce_add3b1_maj3b_wy87;
  assign multm_reduce_add3b1_maj3b_or3b_wx88 = multm_reduce_add3b1_maj3b_wx88 | multm_reduce_add3b1_maj3b_wy88;
  assign multm_reduce_add3b1_maj3b_or3b_wx89 = multm_reduce_add3b1_maj3b_wx89 | multm_reduce_add3b1_maj3b_wy89;
  assign multm_reduce_add3b1_maj3b_or3b_wx90 = multm_reduce_add3b1_maj3b_wx90 | multm_reduce_add3b1_maj3b_wy90;
  assign multm_reduce_add3b1_maj3b_or3b_wx91 = multm_reduce_add3b1_maj3b_wx91 | multm_reduce_add3b1_maj3b_wy91;
  assign multm_reduce_add3b1_maj3b_or3b_wx92 = multm_reduce_add3b1_maj3b_wx92 | multm_reduce_add3b1_maj3b_wy92;
  assign multm_reduce_add3b1_maj3b_or3b_wx93 = multm_reduce_add3b1_maj3b_wx93 | multm_reduce_add3b1_maj3b_wy93;
  assign multm_reduce_add3b1_maj3b_or3b_wx94 = multm_reduce_add3b1_maj3b_wx94 | multm_reduce_add3b1_maj3b_wy94;
  assign multm_reduce_add3b1_maj3b_or3b_wx95 = multm_reduce_add3b1_maj3b_wx95 | multm_reduce_add3b1_maj3b_wy95;
  assign multm_reduce_add3b1_maj3b_or3b_wx96 = multm_reduce_add3b1_maj3b_wx96 | multm_reduce_add3b1_maj3b_wy96;
  assign multm_reduce_add3b1_maj3b_or3b_wx97 = multm_reduce_add3b1_maj3b_wx97 | multm_reduce_add3b1_maj3b_wy97;
  assign multm_reduce_add3b1_maj3b_or3b_wx98 = multm_reduce_add3b1_maj3b_wx98 | multm_reduce_add3b1_maj3b_wy98;
  assign multm_reduce_add3b1_maj3b_or3b_wx99 = multm_reduce_add3b1_maj3b_wx99 | multm_reduce_add3b1_maj3b_wy99;
  assign multm_reduce_add3b1_maj3b_or3b_wx100 = multm_reduce_add3b1_maj3b_wx100 | multm_reduce_add3b1_maj3b_wy100;
  assign multm_reduce_add3b1_maj3b_or3b_wx101 = multm_reduce_add3b1_maj3b_wx101 | multm_reduce_add3b1_maj3b_wy101;
  assign multm_reduce_add3b1_maj3b_or3b_wx102 = multm_reduce_add3b1_maj3b_wx102 | multm_reduce_add3b1_maj3b_wy102;
  assign multm_reduce_add3b1_maj3b_or3b_wx103 = multm_reduce_add3b1_maj3b_wx103 | multm_reduce_add3b1_maj3b_wy103;
  assign multm_reduce_add3b1_maj3b_or3b_wx104 = multm_reduce_add3b1_maj3b_wx104 | multm_reduce_add3b1_maj3b_wy104;
  assign multm_reduce_add3b1_maj3b_or3b_wx105 = multm_reduce_add3b1_maj3b_wx105 | multm_reduce_add3b1_maj3b_wy105;
  assign multm_reduce_add3b1_maj3b_or3b_wx106 = multm_reduce_add3b1_maj3b_wx106 | multm_reduce_add3b1_maj3b_wy106;
  assign multm_reduce_add3b1_maj3b_or3b_wx107 = multm_reduce_add3b1_maj3b_wx107 | multm_reduce_add3b1_maj3b_wy107;
  assign multm_reduce_add3b1_maj3b_or3b_wx108 = multm_reduce_add3b1_maj3b_wx108 | multm_reduce_add3b1_maj3b_wy108;
  assign multm_reduce_add3b1_maj3b_or3b_wx109 = multm_reduce_add3b1_maj3b_wx109 | multm_reduce_add3b1_maj3b_wy109;
  assign multm_reduce_add3b1_maj3b_or3b_wx110 = multm_reduce_add3b1_maj3b_wx110 | multm_reduce_add3b1_maj3b_wy110;
  assign multm_reduce_add3b1_maj3b_or3b_wx111 = multm_reduce_add3b1_maj3b_wx111 | multm_reduce_add3b1_maj3b_wy111;
  assign multm_reduce_add3b1_maj3b_or3b_wx112 = multm_reduce_add3b1_maj3b_wx112 | multm_reduce_add3b1_maj3b_wy112;
  assign multm_reduce_add3b1_maj3b_or3b_wx113 = multm_reduce_add3b1_maj3b_wx113 | multm_reduce_add3b1_maj3b_wy113;
  assign multm_reduce_add3b1_maj3b_or3b_wx114 = multm_reduce_add3b1_maj3b_wx114 | multm_reduce_add3b1_maj3b_wy114;
  assign multm_reduce_add3b1_maj3b_or3b_wx115 = multm_reduce_add3b1_maj3b_wx115 | multm_reduce_add3b1_maj3b_wy115;
  assign multm_reduce_add3b1_maj3b_or3b_wx116 = multm_reduce_add3b1_maj3b_wx116 | multm_reduce_add3b1_maj3b_wy116;
  assign multm_reduce_add3b1_maj3b_or3b_wx117 = multm_reduce_add3b1_maj3b_wx117 | multm_reduce_add3b1_maj3b_wy117;
  assign multm_reduce_add3b1_maj3b_or3b_wx118 = multm_reduce_add3b1_maj3b_wx118 | multm_reduce_add3b1_maj3b_wy118;
  assign multm_reduce_add3b1_maj3b_or3b_wx119 = multm_reduce_add3b1_maj3b_wx119 | multm_reduce_add3b1_maj3b_wy119;
  assign multm_reduce_add3b1_maj3b_or3b_wx120 = multm_reduce_add3b1_maj3b_wx120 | multm_reduce_add3b1_maj3b_wy120;
  assign multm_reduce_add3b1_maj3b_or3b_wx121 = multm_reduce_add3b1_maj3b_wx121 | multm_reduce_add3b1_maj3b_wy121;
  assign multm_reduce_add3b1_maj3b_or3b_wx122 = multm_reduce_add3b1_maj3b_wx122 | multm_reduce_add3b1_maj3b_wy122;
  assign multm_reduce_add3b1_maj3b_or3b_wx123 = multm_reduce_add3b1_maj3b_wx123 | multm_reduce_add3b1_maj3b_wy123;
  assign multm_reduce_add3b1_maj3b_or3b_wx124 = multm_reduce_add3b1_maj3b_wx124 | multm_reduce_add3b1_maj3b_wy124;
  assign multm_reduce_add3b1_maj3b_or3b_wx125 = multm_reduce_add3b1_maj3b_wx125 | multm_reduce_add3b1_maj3b_wy125;
  assign multm_reduce_add3b1_maj3b_or3b_wx126 = multm_reduce_add3b1_maj3b_wx126 | multm_reduce_add3b1_maj3b_wy126;
  assign multm_reduce_add3b1_maj3b_or3b_wx127 = multm_reduce_add3b1_maj3b_wx127 | multm_reduce_add3b1_maj3b_wy127;
  assign multm_reduce_add3b1_maj3b_or3b_wx128 = multm_reduce_add3b1_maj3b_wx128 | multm_reduce_add3b1_maj3b_wy128;
  assign multm_reduce_add3b1_maj3b_or3b_wx129 = multm_reduce_add3b1_maj3b_wx129 | multm_reduce_add3b1_maj3b_wy129;
  assign multm_reduce_add3b1_maj3b_or3b_wx130 = multm_reduce_add3b1_maj3b_wx130 | multm_reduce_add3b1_maj3b_wy130;
  assign multm_reduce_add3b1_maj3b_or3b_wx131 = multm_reduce_add3b1_maj3b_wx131 | multm_reduce_add3b1_maj3b_wy131;
  assign multm_reduce_add3b1_maj3b_or3b_wx132 = multm_reduce_add3b1_maj3b_wx132 | multm_reduce_add3b1_maj3b_wy132;
  assign multm_reduce_add3b1_maj3b_or3b_wx133 = multm_reduce_add3b1_maj3b_wx133 | multm_reduce_add3b1_maj3b_wy133;
  assign multm_reduce_add3b1_maj3b_or3b_wx134 = multm_reduce_add3b1_maj3b_wx134 | multm_reduce_add3b1_maj3b_wy134;
  assign multm_reduce_add3b1_maj3b_or3b_wx135 = multm_reduce_add3b1_maj3b_wx135 | multm_reduce_add3b1_maj3b_wy135;
  assign multm_reduce_add3b1_maj3b_or3b_wx136 = multm_reduce_add3b1_maj3b_wx136 | multm_reduce_add3b1_maj3b_wy136;
  assign multm_reduce_add3b1_maj3b_or3b_wx137 = multm_reduce_add3b1_maj3b_wx137 | multm_reduce_add3b1_maj3b_wy137;
  assign multm_reduce_add3b1_maj3b_or3b_wx138 = multm_reduce_add3b1_maj3b_wx138 | multm_reduce_add3b1_maj3b_wy138;
  assign multm_reduce_add3b1_maj3b_or3b_wx139 = multm_reduce_add3b1_maj3b_wx139 | multm_reduce_add3b1_maj3b_wy139;
  assign multm_reduce_add3b1_maj3b_or3b_wx140 = multm_reduce_add3b1_maj3b_wx140 | multm_reduce_add3b1_maj3b_wy140;
  assign multm_reduce_add3b1_maj3b_or3b_wx141 = multm_reduce_add3b1_maj3b_wx141 | multm_reduce_add3b1_maj3b_wy141;
  assign multm_reduce_add3b1_maj3b_or3b_wx142 = multm_reduce_add3b1_maj3b_wx142 | multm_reduce_add3b1_maj3b_wy142;
  assign multm_reduce_add3b1_maj3b_or3b_wx143 = multm_reduce_add3b1_maj3b_wx143 | multm_reduce_add3b1_maj3b_wy143;
  assign multm_reduce_add3b1_maj3b_or3b_wx144 = multm_reduce_add3b1_maj3b_wx144 | multm_reduce_add3b1_maj3b_wy144;
  assign multm_reduce_add3b1_maj3b_or3b_wx145 = multm_reduce_add3b1_maj3b_wx145 | multm_reduce_add3b1_maj3b_wy145;
  assign multm_reduce_add3b1_maj3b_or3b_wx146 = multm_reduce_add3b1_maj3b_wx146 | multm_reduce_add3b1_maj3b_wy146;
  assign multm_reduce_add3b1_maj3b_or3b_wx147 = multm_reduce_add3b1_maj3b_wx147 | multm_reduce_add3b1_maj3b_wy147;
  assign multm_reduce_add3b1_maj3b_or3b_wx148 = multm_reduce_add3b1_maj3b_wx148 | multm_reduce_add3b1_maj3b_wy148;
  assign multm_reduce_add3b1_maj3b_or3b_wx149 = multm_reduce_add3b1_maj3b_wx149 | multm_reduce_add3b1_maj3b_wy149;
  assign multm_reduce_add3b1_maj3b_or3b_wx150 = multm_reduce_add3b1_maj3b_wx150 | multm_reduce_add3b1_maj3b_wy150;
  assign multm_reduce_add3b1_maj3b_or3b_wx151 = multm_reduce_add3b1_maj3b_wx151 | multm_reduce_add3b1_maj3b_wy151;
  assign multm_reduce_add3b1_maj3b_or3b_wx152 = multm_reduce_add3b1_maj3b_wx152 | multm_reduce_add3b1_maj3b_wy152;
  assign multm_reduce_add3b1_maj3b_or3b_wx153 = multm_reduce_add3b1_maj3b_wx153 | multm_reduce_add3b1_maj3b_wy153;
  assign multm_reduce_add3b1_maj3b_or3b_wx154 = multm_reduce_add3b1_maj3b_wx154 | multm_reduce_add3b1_maj3b_wy154;
  assign multm_reduce_add3b1_maj3b_or3b_wx155 = multm_reduce_add3b1_maj3b_wx155 | multm_reduce_add3b1_maj3b_wy155;
  assign multm_reduce_add3b1_maj3b_or3b_wx156 = multm_reduce_add3b1_maj3b_wx156 | multm_reduce_add3b1_maj3b_wy156;
  assign multm_reduce_add3b1_maj3b_or3b_wx157 = multm_reduce_add3b1_maj3b_wx157 | multm_reduce_add3b1_maj3b_wy157;
  assign multm_reduce_add3b1_maj3b_or3b_wx158 = multm_reduce_add3b1_maj3b_wx158 | multm_reduce_add3b1_maj3b_wy158;
  assign multm_reduce_add3b1_maj3b_or3b_wx159 = multm_reduce_add3b1_maj3b_wx159 | multm_reduce_add3b1_maj3b_wy159;
  assign multm_reduce_add3b1_maj3b_or3b_wx160 = multm_reduce_add3b1_maj3b_wx160 | multm_reduce_add3b1_maj3b_wy160;
  assign multm_reduce_add3b1_maj3b_or3b_wx161 = multm_reduce_add3b1_maj3b_wx161 | multm_reduce_add3b1_maj3b_wy161;
  assign multm_reduce_add3b1_maj3b_or3b_wx162 = multm_reduce_add3b1_maj3b_wx162 | multm_reduce_add3b1_maj3b_wy162;
  assign multm_reduce_add3b1_maj3b_or3b_wx163 = multm_reduce_add3b1_maj3b_wx163 | multm_reduce_add3b1_maj3b_wy163;
  assign multm_reduce_add3b1_maj3b_or3b_wx164 = multm_reduce_add3b1_maj3b_wx164 | multm_reduce_add3b1_maj3b_wy164;
  assign multm_reduce_add3b1_maj3b_or3b_wx165 = multm_reduce_add3b1_maj3b_wx165 | multm_reduce_add3b1_maj3b_wy165;
  assign multm_reduce_add3b1_maj3b_or3b_wx166 = multm_reduce_add3b1_maj3b_wx166 | multm_reduce_add3b1_maj3b_wy166;
  assign multm_reduce_add3b1_maj3b_or3b_wx167 = multm_reduce_add3b1_maj3b_wx167 | multm_reduce_add3b1_maj3b_wy167;
  assign multm_reduce_add3b1_maj3b_or3b_wx168 = multm_reduce_add3b1_maj3b_wx168 | multm_reduce_add3b1_maj3b_wy168;
  assign multm_reduce_add3b1_maj3b_or3b_wx169 = multm_reduce_add3b1_maj3b_wx169 | multm_reduce_add3b1_maj3b_wy169;
  assign multm_reduce_add3b1_maj3b_or3b_wx170 = multm_reduce_add3b1_maj3b_wx170 | multm_reduce_add3b1_maj3b_wy170;
  assign multm_reduce_add3b1_maj3b_or3b_wx171 = multm_reduce_add3b1_maj3b_wx171 | multm_reduce_add3b1_maj3b_wy171;
  assign multm_reduce_add3b1_maj3b_or3b_wx172 = multm_reduce_add3b1_maj3b_wx172 | multm_reduce_add3b1_maj3b_wy172;
  assign multm_reduce_add3b1_maj3b_wx0 = multm_reduce_sb0 & multm_reduce_ms11;
  assign multm_reduce_add3b1_maj3b_wx1 = multm_reduce_sb1 & multm_reduce_ms12;
  assign multm_reduce_add3b1_maj3b_wx2 = multm_reduce_sb2 & multm_reduce_ms13;
  assign multm_reduce_add3b1_maj3b_wx3 = multm_reduce_sb3 & multm_reduce_ms14;
  assign multm_reduce_add3b1_maj3b_wx4 = multm_reduce_sb4 & multm_reduce_ms15;
  assign multm_reduce_add3b1_maj3b_wx5 = multm_reduce_sb5 & multm_reduce_ms16;
  assign multm_reduce_add3b1_maj3b_wx6 = multm_reduce_sb6 & multm_reduce_ms17;
  assign multm_reduce_add3b1_maj3b_wx7 = multm_reduce_sb7 & multm_reduce_ms18;
  assign multm_reduce_add3b1_maj3b_wx8 = multm_reduce_sb8 & multm_reduce_ms19;
  assign multm_reduce_add3b1_maj3b_wx9 = multm_reduce_sb9 & multm_reduce_ms20;
  assign multm_reduce_add3b1_maj3b_wx10 = multm_reduce_sb10 & multm_reduce_ms21;
  assign multm_reduce_add3b1_maj3b_wx11 = multm_reduce_sb11 & multm_reduce_ms22;
  assign multm_reduce_add3b1_maj3b_wx12 = multm_reduce_sb12 & multm_reduce_ms23;
  assign multm_reduce_add3b1_maj3b_wx13 = multm_reduce_sb13 & multm_reduce_ms24;
  assign multm_reduce_add3b1_maj3b_wx14 = multm_reduce_sb14 & multm_reduce_ms25;
  assign multm_reduce_add3b1_maj3b_wx15 = multm_reduce_sb15 & multm_reduce_ms26;
  assign multm_reduce_add3b1_maj3b_wx16 = multm_reduce_sb16 & multm_reduce_ms27;
  assign multm_reduce_add3b1_maj3b_wx17 = multm_reduce_sb17 & multm_reduce_ms28;
  assign multm_reduce_add3b1_maj3b_wx18 = multm_reduce_sb18 & multm_reduce_ms29;
  assign multm_reduce_add3b1_maj3b_wx19 = multm_reduce_sb19 & multm_reduce_ms30;
  assign multm_reduce_add3b1_maj3b_wx20 = multm_reduce_sb20 & multm_reduce_ms31;
  assign multm_reduce_add3b1_maj3b_wx21 = multm_reduce_sb21 & multm_reduce_ms32;
  assign multm_reduce_add3b1_maj3b_wx22 = multm_reduce_sb22 & multm_reduce_ms33;
  assign multm_reduce_add3b1_maj3b_wx23 = multm_reduce_sb23 & multm_reduce_ms34;
  assign multm_reduce_add3b1_maj3b_wx24 = multm_reduce_sb24 & multm_reduce_ms35;
  assign multm_reduce_add3b1_maj3b_wx25 = multm_reduce_sb25 & multm_reduce_ms36;
  assign multm_reduce_add3b1_maj3b_wx26 = multm_reduce_sb26 & multm_reduce_ms37;
  assign multm_reduce_add3b1_maj3b_wx27 = multm_reduce_sb27 & multm_reduce_ms38;
  assign multm_reduce_add3b1_maj3b_wx28 = multm_reduce_sb28 & multm_reduce_ms39;
  assign multm_reduce_add3b1_maj3b_wx29 = multm_reduce_sb29 & multm_reduce_ms40;
  assign multm_reduce_add3b1_maj3b_wx30 = multm_reduce_sb30 & multm_reduce_ms41;
  assign multm_reduce_add3b1_maj3b_wx31 = multm_reduce_sb31 & multm_reduce_ms42;
  assign multm_reduce_add3b1_maj3b_wx32 = multm_reduce_sb32 & multm_reduce_ms43;
  assign multm_reduce_add3b1_maj3b_wx33 = multm_reduce_sb33 & multm_reduce_ms44;
  assign multm_reduce_add3b1_maj3b_wx34 = multm_reduce_sb34 & multm_reduce_ms45;
  assign multm_reduce_add3b1_maj3b_wx35 = multm_reduce_sb35 & multm_reduce_ms46;
  assign multm_reduce_add3b1_maj3b_wx36 = multm_reduce_sb36 & multm_reduce_ms47;
  assign multm_reduce_add3b1_maj3b_wx37 = multm_reduce_sb37 & multm_reduce_ms48;
  assign multm_reduce_add3b1_maj3b_wx38 = multm_reduce_sb38 & multm_reduce_ms49;
  assign multm_reduce_add3b1_maj3b_wx39 = multm_reduce_sb39 & multm_reduce_ms50;
  assign multm_reduce_add3b1_maj3b_wx40 = multm_reduce_sb40 & multm_reduce_ms51;
  assign multm_reduce_add3b1_maj3b_wx41 = multm_reduce_sb41 & multm_reduce_ms52;
  assign multm_reduce_add3b1_maj3b_wx42 = multm_reduce_sb42 & multm_reduce_ms53;
  assign multm_reduce_add3b1_maj3b_wx43 = multm_reduce_sb43 & multm_reduce_ms54;
  assign multm_reduce_add3b1_maj3b_wx44 = multm_reduce_sb44 & multm_reduce_ms55;
  assign multm_reduce_add3b1_maj3b_wx45 = multm_reduce_sb45 & multm_reduce_ms56;
  assign multm_reduce_add3b1_maj3b_wx46 = multm_reduce_sb46 & multm_reduce_ms57;
  assign multm_reduce_add3b1_maj3b_wx47 = multm_reduce_sb47 & multm_reduce_ms58;
  assign multm_reduce_add3b1_maj3b_wx48 = multm_reduce_sb48 & multm_reduce_ms59;
  assign multm_reduce_add3b1_maj3b_wx49 = multm_reduce_sb49 & multm_reduce_ms60;
  assign multm_reduce_add3b1_maj3b_wx50 = multm_reduce_sb50 & multm_reduce_ms61;
  assign multm_reduce_add3b1_maj3b_wx51 = multm_reduce_sb51 & multm_reduce_ms62;
  assign multm_reduce_add3b1_maj3b_wx52 = multm_reduce_sb52 & multm_reduce_ms63;
  assign multm_reduce_add3b1_maj3b_wx53 = multm_reduce_sb53 & multm_reduce_ms64;
  assign multm_reduce_add3b1_maj3b_wx54 = multm_reduce_sb54 & multm_reduce_ms65;
  assign multm_reduce_add3b1_maj3b_wx55 = multm_reduce_sb55 & multm_reduce_ms66;
  assign multm_reduce_add3b1_maj3b_wx56 = multm_reduce_sb56 & multm_reduce_ms67;
  assign multm_reduce_add3b1_maj3b_wx57 = multm_reduce_sb57 & multm_reduce_ms68;
  assign multm_reduce_add3b1_maj3b_wx58 = multm_reduce_sb58 & multm_reduce_ms69;
  assign multm_reduce_add3b1_maj3b_wx59 = multm_reduce_sb59 & multm_reduce_ms70;
  assign multm_reduce_add3b1_maj3b_wx60 = multm_reduce_sb60 & multm_reduce_ms71;
  assign multm_reduce_add3b1_maj3b_wx61 = multm_reduce_sb61 & multm_reduce_ms72;
  assign multm_reduce_add3b1_maj3b_wx62 = multm_reduce_sb62 & multm_reduce_ms73;
  assign multm_reduce_add3b1_maj3b_wx63 = multm_reduce_sb63 & multm_reduce_ms74;
  assign multm_reduce_add3b1_maj3b_wx64 = multm_reduce_sb64 & multm_reduce_ms75;
  assign multm_reduce_add3b1_maj3b_wx65 = multm_reduce_sb65 & multm_reduce_ms76;
  assign multm_reduce_add3b1_maj3b_wx66 = multm_reduce_sb66 & multm_reduce_ms77;
  assign multm_reduce_add3b1_maj3b_wx67 = multm_reduce_sb67 & multm_reduce_ms78;
  assign multm_reduce_add3b1_maj3b_wx68 = multm_reduce_sb68 & multm_reduce_ms79;
  assign multm_reduce_add3b1_maj3b_wx69 = multm_reduce_sb69 & multm_reduce_ms80;
  assign multm_reduce_add3b1_maj3b_wx70 = multm_reduce_sb70 & multm_reduce_ms81;
  assign multm_reduce_add3b1_maj3b_wx71 = multm_reduce_sb71 & multm_reduce_ms82;
  assign multm_reduce_add3b1_maj3b_wx72 = multm_reduce_sb72 & multm_reduce_ms83;
  assign multm_reduce_add3b1_maj3b_wx73 = multm_reduce_sb73 & multm_reduce_ms84;
  assign multm_reduce_add3b1_maj3b_wx74 = multm_reduce_sb74 & multm_reduce_ms85;
  assign multm_reduce_add3b1_maj3b_wx75 = multm_reduce_sb75 & multm_reduce_ms86;
  assign multm_reduce_add3b1_maj3b_wx76 = multm_reduce_sb76 & multm_reduce_ms87;
  assign multm_reduce_add3b1_maj3b_wx77 = multm_reduce_sb77 & multm_reduce_ms88;
  assign multm_reduce_add3b1_maj3b_wx78 = multm_reduce_sb78 & multm_reduce_ms89;
  assign multm_reduce_add3b1_maj3b_wx79 = multm_reduce_sb79 & multm_reduce_ms90;
  assign multm_reduce_add3b1_maj3b_wx80 = multm_reduce_sb80 & multm_reduce_ms91;
  assign multm_reduce_add3b1_maj3b_wx81 = multm_reduce_sb81 & multm_reduce_ms92;
  assign multm_reduce_add3b1_maj3b_wx82 = multm_reduce_sb82 & multm_reduce_ms93;
  assign multm_reduce_add3b1_maj3b_wx83 = multm_reduce_sb83 & multm_reduce_ms94;
  assign multm_reduce_add3b1_maj3b_wx84 = multm_reduce_sb84 & multm_reduce_ms95;
  assign multm_reduce_add3b1_maj3b_wx85 = multm_reduce_sb85 & multm_reduce_ms96;
  assign multm_reduce_add3b1_maj3b_wx86 = multm_reduce_sb86 & multm_reduce_ms97;
  assign multm_reduce_add3b1_maj3b_wx87 = multm_reduce_sb87 & multm_reduce_ms98;
  assign multm_reduce_add3b1_maj3b_wx88 = multm_reduce_sb88 & multm_reduce_ms99;
  assign multm_reduce_add3b1_maj3b_wx89 = multm_reduce_sb89 & multm_reduce_ms100;
  assign multm_reduce_add3b1_maj3b_wx90 = multm_reduce_sb90 & multm_reduce_ms101;
  assign multm_reduce_add3b1_maj3b_wx91 = multm_reduce_sb91 & multm_reduce_ms102;
  assign multm_reduce_add3b1_maj3b_wx92 = multm_reduce_sb92 & multm_reduce_ms103;
  assign multm_reduce_add3b1_maj3b_wx93 = multm_reduce_sb93 & multm_reduce_ms104;
  assign multm_reduce_add3b1_maj3b_wx94 = multm_reduce_sb94 & multm_reduce_ms105;
  assign multm_reduce_add3b1_maj3b_wx95 = multm_reduce_sb95 & multm_reduce_ms106;
  assign multm_reduce_add3b1_maj3b_wx96 = multm_reduce_sb96 & multm_reduce_ms107;
  assign multm_reduce_add3b1_maj3b_wx97 = multm_reduce_sb97 & multm_reduce_ms108;
  assign multm_reduce_add3b1_maj3b_wx98 = multm_reduce_sb98 & multm_reduce_ms109;
  assign multm_reduce_add3b1_maj3b_wx99 = multm_reduce_sb99 & multm_reduce_ms110;
  assign multm_reduce_add3b1_maj3b_wx100 = multm_reduce_sb100 & multm_reduce_ms111;
  assign multm_reduce_add3b1_maj3b_wx101 = multm_reduce_sb101 & multm_reduce_ms112;
  assign multm_reduce_add3b1_maj3b_wx102 = multm_reduce_sb102 & multm_reduce_ms113;
  assign multm_reduce_add3b1_maj3b_wx103 = multm_reduce_sb103 & multm_reduce_ms114;
  assign multm_reduce_add3b1_maj3b_wx104 = multm_reduce_sb104 & multm_reduce_ms115;
  assign multm_reduce_add3b1_maj3b_wx105 = multm_reduce_sb105 & multm_reduce_ms116;
  assign multm_reduce_add3b1_maj3b_wx106 = multm_reduce_sb106 & multm_reduce_ms117;
  assign multm_reduce_add3b1_maj3b_wx107 = multm_reduce_sb107 & multm_reduce_ms118;
  assign multm_reduce_add3b1_maj3b_wx108 = multm_reduce_sb108 & multm_reduce_ms119;
  assign multm_reduce_add3b1_maj3b_wx109 = multm_reduce_sb109 & multm_reduce_ms120;
  assign multm_reduce_add3b1_maj3b_wx110 = multm_reduce_sb110 & multm_reduce_ms121;
  assign multm_reduce_add3b1_maj3b_wx111 = multm_reduce_sb111 & multm_reduce_ms122;
  assign multm_reduce_add3b1_maj3b_wx112 = multm_reduce_sb112 & multm_reduce_ms123;
  assign multm_reduce_add3b1_maj3b_wx113 = multm_reduce_sb113 & multm_reduce_ms124;
  assign multm_reduce_add3b1_maj3b_wx114 = multm_reduce_sb114 & multm_reduce_ms125;
  assign multm_reduce_add3b1_maj3b_wx115 = multm_reduce_sb115 & multm_reduce_ms126;
  assign multm_reduce_add3b1_maj3b_wx116 = multm_reduce_sb116 & multm_reduce_ms127;
  assign multm_reduce_add3b1_maj3b_wx117 = multm_reduce_sb117 & multm_reduce_ms128;
  assign multm_reduce_add3b1_maj3b_wx118 = multm_reduce_sb118 & multm_reduce_ms129;
  assign multm_reduce_add3b1_maj3b_wx119 = multm_reduce_sb119 & multm_reduce_ms130;
  assign multm_reduce_add3b1_maj3b_wx120 = multm_reduce_sb120 & multm_reduce_ms131;
  assign multm_reduce_add3b1_maj3b_wx121 = multm_reduce_sb121 & multm_reduce_ms132;
  assign multm_reduce_add3b1_maj3b_wx122 = multm_reduce_sb122 & multm_reduce_ms133;
  assign multm_reduce_add3b1_maj3b_wx123 = multm_reduce_sb123 & multm_reduce_ms134;
  assign multm_reduce_add3b1_maj3b_wx124 = multm_reduce_sb124 & multm_reduce_ms135;
  assign multm_reduce_add3b1_maj3b_wx125 = multm_reduce_sb125 & multm_reduce_ms136;
  assign multm_reduce_add3b1_maj3b_wx126 = multm_reduce_sb126 & multm_reduce_ms137;
  assign multm_reduce_add3b1_maj3b_wx127 = multm_reduce_sb127 & multm_reduce_ms138;
  assign multm_reduce_add3b1_maj3b_wx128 = multm_reduce_sb128 & multm_reduce_ms139;
  assign multm_reduce_add3b1_maj3b_wx129 = multm_reduce_sb129 & multm_reduce_ms140;
  assign multm_reduce_add3b1_maj3b_wx130 = multm_reduce_sb130 & multm_reduce_ms141;
  assign multm_reduce_add3b1_maj3b_wx131 = multm_reduce_sb131 & multm_reduce_ms142;
  assign multm_reduce_add3b1_maj3b_wx132 = multm_reduce_sb132 & multm_reduce_ms143;
  assign multm_reduce_add3b1_maj3b_wx133 = multm_reduce_sb133 & multm_reduce_ms144;
  assign multm_reduce_add3b1_maj3b_wx134 = multm_reduce_sb134 & multm_reduce_ms145;
  assign multm_reduce_add3b1_maj3b_wx135 = multm_reduce_sb135 & multm_reduce_ms146;
  assign multm_reduce_add3b1_maj3b_wx136 = multm_reduce_sb136 & multm_reduce_ms147;
  assign multm_reduce_add3b1_maj3b_wx137 = multm_reduce_sb137 & multm_reduce_ms148;
  assign multm_reduce_add3b1_maj3b_wx138 = multm_reduce_sb138 & multm_reduce_ms149;
  assign multm_reduce_add3b1_maj3b_wx139 = multm_reduce_sb139 & multm_reduce_ms150;
  assign multm_reduce_add3b1_maj3b_wx140 = multm_reduce_sb140 & multm_reduce_ms151;
  assign multm_reduce_add3b1_maj3b_wx141 = multm_reduce_sb141 & multm_reduce_ms152;
  assign multm_reduce_add3b1_maj3b_wx142 = multm_reduce_sb142 & multm_reduce_ms153;
  assign multm_reduce_add3b1_maj3b_wx143 = multm_reduce_sb143 & multm_reduce_ms154;
  assign multm_reduce_add3b1_maj3b_wx144 = multm_reduce_sb144 & multm_reduce_ms155;
  assign multm_reduce_add3b1_maj3b_wx145 = multm_reduce_sb145 & multm_reduce_ms156;
  assign multm_reduce_add3b1_maj3b_wx146 = multm_reduce_sb146 & multm_reduce_ms157;
  assign multm_reduce_add3b1_maj3b_wx147 = multm_reduce_sb147 & multm_reduce_ms158;
  assign multm_reduce_add3b1_maj3b_wx148 = multm_reduce_sb148 & multm_reduce_ms159;
  assign multm_reduce_add3b1_maj3b_wx149 = multm_reduce_sb149 & multm_reduce_ms160;
  assign multm_reduce_add3b1_maj3b_wx150 = multm_reduce_sb150 & multm_reduce_ms161;
  assign multm_reduce_add3b1_maj3b_wx151 = multm_reduce_sb151 & multm_reduce_ms162;
  assign multm_reduce_add3b1_maj3b_wx152 = multm_reduce_sb152 & multm_reduce_ms163;
  assign multm_reduce_add3b1_maj3b_wx153 = multm_reduce_sb153 & multm_reduce_ms164;
  assign multm_reduce_add3b1_maj3b_wx154 = multm_reduce_sb154 & multm_reduce_ms165;
  assign multm_reduce_add3b1_maj3b_wx155 = multm_reduce_sb155 & multm_reduce_ms166;
  assign multm_reduce_add3b1_maj3b_wx156 = multm_reduce_sb156 & multm_reduce_ms167;
  assign multm_reduce_add3b1_maj3b_wx157 = multm_reduce_sb157 & multm_reduce_ms168;
  assign multm_reduce_add3b1_maj3b_wx158 = multm_reduce_sb158 & multm_reduce_ms169;
  assign multm_reduce_add3b1_maj3b_wx159 = multm_reduce_sb159 & multm_reduce_ms170;
  assign multm_reduce_add3b1_maj3b_wx160 = multm_reduce_sb160 & multm_reduce_ms171;
  assign multm_reduce_add3b1_maj3b_wx161 = multm_reduce_sb161 & multm_reduce_ms172;
  assign multm_reduce_add3b1_maj3b_wx162 = multm_reduce_sb162 & multm_reduce_ms173;
  assign multm_reduce_add3b1_maj3b_wx163 = multm_reduce_sb163 & multm_reduce_ms174;
  assign multm_reduce_add3b1_maj3b_wx164 = multm_reduce_sb164 & multm_reduce_ms175;
  assign multm_reduce_add3b1_maj3b_wx165 = multm_reduce_sb165 & multm_reduce_ms176;
  assign multm_reduce_add3b1_maj3b_wx166 = multm_reduce_sb166 & multm_reduce_ms177;
  assign multm_reduce_add3b1_maj3b_wx167 = multm_reduce_sb167 & multm_reduce_ms178;
  assign multm_reduce_add3b1_maj3b_wx168 = multm_reduce_sb168 & multm_reduce_ms179;
  assign multm_reduce_add3b1_maj3b_wx169 = multm_reduce_sb169 & multm_reduce_ms180;
  assign multm_reduce_add3b1_maj3b_wx170 = multm_reduce_sb170 & multm_reduce_ms181;
  assign multm_reduce_add3b1_maj3b_wx171 = multm_reduce_sb171 & multm_reduce_ms182;
  assign multm_reduce_add3b1_maj3b_wx172 = multm_reduce_sb172 & multm_reduce_ms183;
  assign multm_reduce_add3b1_maj3b_wy0 = multm_reduce_sb0 & multm_reduce_mc10;
  assign multm_reduce_add3b1_maj3b_wy1 = multm_reduce_sb1 & multm_reduce_mc11;
  assign multm_reduce_add3b1_maj3b_wy2 = multm_reduce_sb2 & multm_reduce_mc12;
  assign multm_reduce_add3b1_maj3b_wy3 = multm_reduce_sb3 & multm_reduce_mc13;
  assign multm_reduce_add3b1_maj3b_wy4 = multm_reduce_sb4 & multm_reduce_mc14;
  assign multm_reduce_add3b1_maj3b_wy5 = multm_reduce_sb5 & multm_reduce_mc15;
  assign multm_reduce_add3b1_maj3b_wy6 = multm_reduce_sb6 & multm_reduce_mc16;
  assign multm_reduce_add3b1_maj3b_wy7 = multm_reduce_sb7 & multm_reduce_mc17;
  assign multm_reduce_add3b1_maj3b_wy8 = multm_reduce_sb8 & multm_reduce_mc18;
  assign multm_reduce_add3b1_maj3b_wy9 = multm_reduce_sb9 & multm_reduce_mc19;
  assign multm_reduce_add3b1_maj3b_wy10 = multm_reduce_sb10 & multm_reduce_mc20;
  assign multm_reduce_add3b1_maj3b_wy11 = multm_reduce_sb11 & multm_reduce_mc21;
  assign multm_reduce_add3b1_maj3b_wy12 = multm_reduce_sb12 & multm_reduce_mc22;
  assign multm_reduce_add3b1_maj3b_wy13 = multm_reduce_sb13 & multm_reduce_mc23;
  assign multm_reduce_add3b1_maj3b_wy14 = multm_reduce_sb14 & multm_reduce_mc24;
  assign multm_reduce_add3b1_maj3b_wy15 = multm_reduce_sb15 & multm_reduce_mc25;
  assign multm_reduce_add3b1_maj3b_wy16 = multm_reduce_sb16 & multm_reduce_mc26;
  assign multm_reduce_add3b1_maj3b_wy17 = multm_reduce_sb17 & multm_reduce_mc27;
  assign multm_reduce_add3b1_maj3b_wy18 = multm_reduce_sb18 & multm_reduce_mc28;
  assign multm_reduce_add3b1_maj3b_wy19 = multm_reduce_sb19 & multm_reduce_mc29;
  assign multm_reduce_add3b1_maj3b_wy20 = multm_reduce_sb20 & multm_reduce_mc30;
  assign multm_reduce_add3b1_maj3b_wy21 = multm_reduce_sb21 & multm_reduce_mc31;
  assign multm_reduce_add3b1_maj3b_wy22 = multm_reduce_sb22 & multm_reduce_mc32;
  assign multm_reduce_add3b1_maj3b_wy23 = multm_reduce_sb23 & multm_reduce_mc33;
  assign multm_reduce_add3b1_maj3b_wy24 = multm_reduce_sb24 & multm_reduce_mc34;
  assign multm_reduce_add3b1_maj3b_wy25 = multm_reduce_sb25 & multm_reduce_mc35;
  assign multm_reduce_add3b1_maj3b_wy26 = multm_reduce_sb26 & multm_reduce_mc36;
  assign multm_reduce_add3b1_maj3b_wy27 = multm_reduce_sb27 & multm_reduce_mc37;
  assign multm_reduce_add3b1_maj3b_wy28 = multm_reduce_sb28 & multm_reduce_mc38;
  assign multm_reduce_add3b1_maj3b_wy29 = multm_reduce_sb29 & multm_reduce_mc39;
  assign multm_reduce_add3b1_maj3b_wy30 = multm_reduce_sb30 & multm_reduce_mc40;
  assign multm_reduce_add3b1_maj3b_wy31 = multm_reduce_sb31 & multm_reduce_mc41;
  assign multm_reduce_add3b1_maj3b_wy32 = multm_reduce_sb32 & multm_reduce_mc42;
  assign multm_reduce_add3b1_maj3b_wy33 = multm_reduce_sb33 & multm_reduce_mc43;
  assign multm_reduce_add3b1_maj3b_wy34 = multm_reduce_sb34 & multm_reduce_mc44;
  assign multm_reduce_add3b1_maj3b_wy35 = multm_reduce_sb35 & multm_reduce_mc45;
  assign multm_reduce_add3b1_maj3b_wy36 = multm_reduce_sb36 & multm_reduce_mc46;
  assign multm_reduce_add3b1_maj3b_wy37 = multm_reduce_sb37 & multm_reduce_mc47;
  assign multm_reduce_add3b1_maj3b_wy38 = multm_reduce_sb38 & multm_reduce_mc48;
  assign multm_reduce_add3b1_maj3b_wy39 = multm_reduce_sb39 & multm_reduce_mc49;
  assign multm_reduce_add3b1_maj3b_wy40 = multm_reduce_sb40 & multm_reduce_mc50;
  assign multm_reduce_add3b1_maj3b_wy41 = multm_reduce_sb41 & multm_reduce_mc51;
  assign multm_reduce_add3b1_maj3b_wy42 = multm_reduce_sb42 & multm_reduce_mc52;
  assign multm_reduce_add3b1_maj3b_wy43 = multm_reduce_sb43 & multm_reduce_mc53;
  assign multm_reduce_add3b1_maj3b_wy44 = multm_reduce_sb44 & multm_reduce_mc54;
  assign multm_reduce_add3b1_maj3b_wy45 = multm_reduce_sb45 & multm_reduce_mc55;
  assign multm_reduce_add3b1_maj3b_wy46 = multm_reduce_sb46 & multm_reduce_mc56;
  assign multm_reduce_add3b1_maj3b_wy47 = multm_reduce_sb47 & multm_reduce_mc57;
  assign multm_reduce_add3b1_maj3b_wy48 = multm_reduce_sb48 & multm_reduce_mc58;
  assign multm_reduce_add3b1_maj3b_wy49 = multm_reduce_sb49 & multm_reduce_mc59;
  assign multm_reduce_add3b1_maj3b_wy50 = multm_reduce_sb50 & multm_reduce_mc60;
  assign multm_reduce_add3b1_maj3b_wy51 = multm_reduce_sb51 & multm_reduce_mc61;
  assign multm_reduce_add3b1_maj3b_wy52 = multm_reduce_sb52 & multm_reduce_mc62;
  assign multm_reduce_add3b1_maj3b_wy53 = multm_reduce_sb53 & multm_reduce_mc63;
  assign multm_reduce_add3b1_maj3b_wy54 = multm_reduce_sb54 & multm_reduce_mc64;
  assign multm_reduce_add3b1_maj3b_wy55 = multm_reduce_sb55 & multm_reduce_mc65;
  assign multm_reduce_add3b1_maj3b_wy56 = multm_reduce_sb56 & multm_reduce_mc66;
  assign multm_reduce_add3b1_maj3b_wy57 = multm_reduce_sb57 & multm_reduce_mc67;
  assign multm_reduce_add3b1_maj3b_wy58 = multm_reduce_sb58 & multm_reduce_mc68;
  assign multm_reduce_add3b1_maj3b_wy59 = multm_reduce_sb59 & multm_reduce_mc69;
  assign multm_reduce_add3b1_maj3b_wy60 = multm_reduce_sb60 & multm_reduce_mc70;
  assign multm_reduce_add3b1_maj3b_wy61 = multm_reduce_sb61 & multm_reduce_mc71;
  assign multm_reduce_add3b1_maj3b_wy62 = multm_reduce_sb62 & multm_reduce_mc72;
  assign multm_reduce_add3b1_maj3b_wy63 = multm_reduce_sb63 & multm_reduce_mc73;
  assign multm_reduce_add3b1_maj3b_wy64 = multm_reduce_sb64 & multm_reduce_mc74;
  assign multm_reduce_add3b1_maj3b_wy65 = multm_reduce_sb65 & multm_reduce_mc75;
  assign multm_reduce_add3b1_maj3b_wy66 = multm_reduce_sb66 & multm_reduce_mc76;
  assign multm_reduce_add3b1_maj3b_wy67 = multm_reduce_sb67 & multm_reduce_mc77;
  assign multm_reduce_add3b1_maj3b_wy68 = multm_reduce_sb68 & multm_reduce_mc78;
  assign multm_reduce_add3b1_maj3b_wy69 = multm_reduce_sb69 & multm_reduce_mc79;
  assign multm_reduce_add3b1_maj3b_wy70 = multm_reduce_sb70 & multm_reduce_mc80;
  assign multm_reduce_add3b1_maj3b_wy71 = multm_reduce_sb71 & multm_reduce_mc81;
  assign multm_reduce_add3b1_maj3b_wy72 = multm_reduce_sb72 & multm_reduce_mc82;
  assign multm_reduce_add3b1_maj3b_wy73 = multm_reduce_sb73 & multm_reduce_mc83;
  assign multm_reduce_add3b1_maj3b_wy74 = multm_reduce_sb74 & multm_reduce_mc84;
  assign multm_reduce_add3b1_maj3b_wy75 = multm_reduce_sb75 & multm_reduce_mc85;
  assign multm_reduce_add3b1_maj3b_wy76 = multm_reduce_sb76 & multm_reduce_mc86;
  assign multm_reduce_add3b1_maj3b_wy77 = multm_reduce_sb77 & multm_reduce_mc87;
  assign multm_reduce_add3b1_maj3b_wy78 = multm_reduce_sb78 & multm_reduce_mc88;
  assign multm_reduce_add3b1_maj3b_wy79 = multm_reduce_sb79 & multm_reduce_mc89;
  assign multm_reduce_add3b1_maj3b_wy80 = multm_reduce_sb80 & multm_reduce_mc90;
  assign multm_reduce_add3b1_maj3b_wy81 = multm_reduce_sb81 & multm_reduce_mc91;
  assign multm_reduce_add3b1_maj3b_wy82 = multm_reduce_sb82 & multm_reduce_mc92;
  assign multm_reduce_add3b1_maj3b_wy83 = multm_reduce_sb83 & multm_reduce_mc93;
  assign multm_reduce_add3b1_maj3b_wy84 = multm_reduce_sb84 & multm_reduce_mc94;
  assign multm_reduce_add3b1_maj3b_wy85 = multm_reduce_sb85 & multm_reduce_mc95;
  assign multm_reduce_add3b1_maj3b_wy86 = multm_reduce_sb86 & multm_reduce_mc96;
  assign multm_reduce_add3b1_maj3b_wy87 = multm_reduce_sb87 & multm_reduce_mc97;
  assign multm_reduce_add3b1_maj3b_wy88 = multm_reduce_sb88 & multm_reduce_mc98;
  assign multm_reduce_add3b1_maj3b_wy89 = multm_reduce_sb89 & multm_reduce_mc99;
  assign multm_reduce_add3b1_maj3b_wy90 = multm_reduce_sb90 & multm_reduce_mc100;
  assign multm_reduce_add3b1_maj3b_wy91 = multm_reduce_sb91 & multm_reduce_mc101;
  assign multm_reduce_add3b1_maj3b_wy92 = multm_reduce_sb92 & multm_reduce_mc102;
  assign multm_reduce_add3b1_maj3b_wy93 = multm_reduce_sb93 & multm_reduce_mc103;
  assign multm_reduce_add3b1_maj3b_wy94 = multm_reduce_sb94 & multm_reduce_mc104;
  assign multm_reduce_add3b1_maj3b_wy95 = multm_reduce_sb95 & multm_reduce_mc105;
  assign multm_reduce_add3b1_maj3b_wy96 = multm_reduce_sb96 & multm_reduce_mc106;
  assign multm_reduce_add3b1_maj3b_wy97 = multm_reduce_sb97 & multm_reduce_mc107;
  assign multm_reduce_add3b1_maj3b_wy98 = multm_reduce_sb98 & multm_reduce_mc108;
  assign multm_reduce_add3b1_maj3b_wy99 = multm_reduce_sb99 & multm_reduce_mc109;
  assign multm_reduce_add3b1_maj3b_wy100 = multm_reduce_sb100 & multm_reduce_mc110;
  assign multm_reduce_add3b1_maj3b_wy101 = multm_reduce_sb101 & multm_reduce_mc111;
  assign multm_reduce_add3b1_maj3b_wy102 = multm_reduce_sb102 & multm_reduce_mc112;
  assign multm_reduce_add3b1_maj3b_wy103 = multm_reduce_sb103 & multm_reduce_mc113;
  assign multm_reduce_add3b1_maj3b_wy104 = multm_reduce_sb104 & multm_reduce_mc114;
  assign multm_reduce_add3b1_maj3b_wy105 = multm_reduce_sb105 & multm_reduce_mc115;
  assign multm_reduce_add3b1_maj3b_wy106 = multm_reduce_sb106 & multm_reduce_mc116;
  assign multm_reduce_add3b1_maj3b_wy107 = multm_reduce_sb107 & multm_reduce_mc117;
  assign multm_reduce_add3b1_maj3b_wy108 = multm_reduce_sb108 & multm_reduce_mc118;
  assign multm_reduce_add3b1_maj3b_wy109 = multm_reduce_sb109 & multm_reduce_mc119;
  assign multm_reduce_add3b1_maj3b_wy110 = multm_reduce_sb110 & multm_reduce_mc120;
  assign multm_reduce_add3b1_maj3b_wy111 = multm_reduce_sb111 & multm_reduce_mc121;
  assign multm_reduce_add3b1_maj3b_wy112 = multm_reduce_sb112 & multm_reduce_mc122;
  assign multm_reduce_add3b1_maj3b_wy113 = multm_reduce_sb113 & multm_reduce_mc123;
  assign multm_reduce_add3b1_maj3b_wy114 = multm_reduce_sb114 & multm_reduce_mc124;
  assign multm_reduce_add3b1_maj3b_wy115 = multm_reduce_sb115 & multm_reduce_mc125;
  assign multm_reduce_add3b1_maj3b_wy116 = multm_reduce_sb116 & multm_reduce_mc126;
  assign multm_reduce_add3b1_maj3b_wy117 = multm_reduce_sb117 & multm_reduce_mc127;
  assign multm_reduce_add3b1_maj3b_wy118 = multm_reduce_sb118 & multm_reduce_mc128;
  assign multm_reduce_add3b1_maj3b_wy119 = multm_reduce_sb119 & multm_reduce_mc129;
  assign multm_reduce_add3b1_maj3b_wy120 = multm_reduce_sb120 & multm_reduce_mc130;
  assign multm_reduce_add3b1_maj3b_wy121 = multm_reduce_sb121 & multm_reduce_mc131;
  assign multm_reduce_add3b1_maj3b_wy122 = multm_reduce_sb122 & multm_reduce_mc132;
  assign multm_reduce_add3b1_maj3b_wy123 = multm_reduce_sb123 & multm_reduce_mc133;
  assign multm_reduce_add3b1_maj3b_wy124 = multm_reduce_sb124 & multm_reduce_mc134;
  assign multm_reduce_add3b1_maj3b_wy125 = multm_reduce_sb125 & multm_reduce_mc135;
  assign multm_reduce_add3b1_maj3b_wy126 = multm_reduce_sb126 & multm_reduce_mc136;
  assign multm_reduce_add3b1_maj3b_wy127 = multm_reduce_sb127 & multm_reduce_mc137;
  assign multm_reduce_add3b1_maj3b_wy128 = multm_reduce_sb128 & multm_reduce_mc138;
  assign multm_reduce_add3b1_maj3b_wy129 = multm_reduce_sb129 & multm_reduce_mc139;
  assign multm_reduce_add3b1_maj3b_wy130 = multm_reduce_sb130 & multm_reduce_mc140;
  assign multm_reduce_add3b1_maj3b_wy131 = multm_reduce_sb131 & multm_reduce_mc141;
  assign multm_reduce_add3b1_maj3b_wy132 = multm_reduce_sb132 & multm_reduce_mc142;
  assign multm_reduce_add3b1_maj3b_wy133 = multm_reduce_sb133 & multm_reduce_mc143;
  assign multm_reduce_add3b1_maj3b_wy134 = multm_reduce_sb134 & multm_reduce_mc144;
  assign multm_reduce_add3b1_maj3b_wy135 = multm_reduce_sb135 & multm_reduce_mc145;
  assign multm_reduce_add3b1_maj3b_wy136 = multm_reduce_sb136 & multm_reduce_mc146;
  assign multm_reduce_add3b1_maj3b_wy137 = multm_reduce_sb137 & multm_reduce_mc147;
  assign multm_reduce_add3b1_maj3b_wy138 = multm_reduce_sb138 & multm_reduce_mc148;
  assign multm_reduce_add3b1_maj3b_wy139 = multm_reduce_sb139 & multm_reduce_mc149;
  assign multm_reduce_add3b1_maj3b_wy140 = multm_reduce_sb140 & multm_reduce_mc150;
  assign multm_reduce_add3b1_maj3b_wy141 = multm_reduce_sb141 & multm_reduce_mc151;
  assign multm_reduce_add3b1_maj3b_wy142 = multm_reduce_sb142 & multm_reduce_mc152;
  assign multm_reduce_add3b1_maj3b_wy143 = multm_reduce_sb143 & multm_reduce_mc153;
  assign multm_reduce_add3b1_maj3b_wy144 = multm_reduce_sb144 & multm_reduce_mc154;
  assign multm_reduce_add3b1_maj3b_wy145 = multm_reduce_sb145 & multm_reduce_mc155;
  assign multm_reduce_add3b1_maj3b_wy146 = multm_reduce_sb146 & multm_reduce_mc156;
  assign multm_reduce_add3b1_maj3b_wy147 = multm_reduce_sb147 & multm_reduce_mc157;
  assign multm_reduce_add3b1_maj3b_wy148 = multm_reduce_sb148 & multm_reduce_mc158;
  assign multm_reduce_add3b1_maj3b_wy149 = multm_reduce_sb149 & multm_reduce_mc159;
  assign multm_reduce_add3b1_maj3b_wy150 = multm_reduce_sb150 & multm_reduce_mc160;
  assign multm_reduce_add3b1_maj3b_wy151 = multm_reduce_sb151 & multm_reduce_mc161;
  assign multm_reduce_add3b1_maj3b_wy152 = multm_reduce_sb152 & multm_reduce_mc162;
  assign multm_reduce_add3b1_maj3b_wy153 = multm_reduce_sb153 & multm_reduce_mc163;
  assign multm_reduce_add3b1_maj3b_wy154 = multm_reduce_sb154 & multm_reduce_mc164;
  assign multm_reduce_add3b1_maj3b_wy155 = multm_reduce_sb155 & multm_reduce_mc165;
  assign multm_reduce_add3b1_maj3b_wy156 = multm_reduce_sb156 & multm_reduce_mc166;
  assign multm_reduce_add3b1_maj3b_wy157 = multm_reduce_sb157 & multm_reduce_mc167;
  assign multm_reduce_add3b1_maj3b_wy158 = multm_reduce_sb158 & multm_reduce_mc168;
  assign multm_reduce_add3b1_maj3b_wy159 = multm_reduce_sb159 & multm_reduce_mc169;
  assign multm_reduce_add3b1_maj3b_wy160 = multm_reduce_sb160 & multm_reduce_mc170;
  assign multm_reduce_add3b1_maj3b_wy161 = multm_reduce_sb161 & multm_reduce_mc171;
  assign multm_reduce_add3b1_maj3b_wy162 = multm_reduce_sb162 & multm_reduce_mc172;
  assign multm_reduce_add3b1_maj3b_wy163 = multm_reduce_sb163 & multm_reduce_mc173;
  assign multm_reduce_add3b1_maj3b_wy164 = multm_reduce_sb164 & multm_reduce_mc174;
  assign multm_reduce_add3b1_maj3b_wy165 = multm_reduce_sb165 & multm_reduce_mc175;
  assign multm_reduce_add3b1_maj3b_wy166 = multm_reduce_sb166 & multm_reduce_mc176;
  assign multm_reduce_add3b1_maj3b_wy167 = multm_reduce_sb167 & multm_reduce_mc177;
  assign multm_reduce_add3b1_maj3b_wy168 = multm_reduce_sb168 & multm_reduce_mc178;
  assign multm_reduce_add3b1_maj3b_wy169 = multm_reduce_sb169 & multm_reduce_mc179;
  assign multm_reduce_add3b1_maj3b_wy170 = multm_reduce_sb170 & multm_reduce_mc180;
  assign multm_reduce_add3b1_maj3b_wy171 = multm_reduce_sb171 & multm_reduce_mc181;
  assign multm_reduce_add3b1_maj3b_wy172 = multm_reduce_sb172 & multm_reduce_mc182;
  assign multm_reduce_add3b1_maj3b_xy0 = multm_reduce_ms11 & multm_reduce_mc10;
  assign multm_reduce_add3b1_maj3b_xy1 = multm_reduce_ms12 & multm_reduce_mc11;
  assign multm_reduce_add3b1_maj3b_xy2 = multm_reduce_ms13 & multm_reduce_mc12;
  assign multm_reduce_add3b1_maj3b_xy3 = multm_reduce_ms14 & multm_reduce_mc13;
  assign multm_reduce_add3b1_maj3b_xy4 = multm_reduce_ms15 & multm_reduce_mc14;
  assign multm_reduce_add3b1_maj3b_xy5 = multm_reduce_ms16 & multm_reduce_mc15;
  assign multm_reduce_add3b1_maj3b_xy6 = multm_reduce_ms17 & multm_reduce_mc16;
  assign multm_reduce_add3b1_maj3b_xy7 = multm_reduce_ms18 & multm_reduce_mc17;
  assign multm_reduce_add3b1_maj3b_xy8 = multm_reduce_ms19 & multm_reduce_mc18;
  assign multm_reduce_add3b1_maj3b_xy9 = multm_reduce_ms20 & multm_reduce_mc19;
  assign multm_reduce_add3b1_maj3b_xy10 = multm_reduce_ms21 & multm_reduce_mc20;
  assign multm_reduce_add3b1_maj3b_xy11 = multm_reduce_ms22 & multm_reduce_mc21;
  assign multm_reduce_add3b1_maj3b_xy12 = multm_reduce_ms23 & multm_reduce_mc22;
  assign multm_reduce_add3b1_maj3b_xy13 = multm_reduce_ms24 & multm_reduce_mc23;
  assign multm_reduce_add3b1_maj3b_xy14 = multm_reduce_ms25 & multm_reduce_mc24;
  assign multm_reduce_add3b1_maj3b_xy15 = multm_reduce_ms26 & multm_reduce_mc25;
  assign multm_reduce_add3b1_maj3b_xy16 = multm_reduce_ms27 & multm_reduce_mc26;
  assign multm_reduce_add3b1_maj3b_xy17 = multm_reduce_ms28 & multm_reduce_mc27;
  assign multm_reduce_add3b1_maj3b_xy18 = multm_reduce_ms29 & multm_reduce_mc28;
  assign multm_reduce_add3b1_maj3b_xy19 = multm_reduce_ms30 & multm_reduce_mc29;
  assign multm_reduce_add3b1_maj3b_xy20 = multm_reduce_ms31 & multm_reduce_mc30;
  assign multm_reduce_add3b1_maj3b_xy21 = multm_reduce_ms32 & multm_reduce_mc31;
  assign multm_reduce_add3b1_maj3b_xy22 = multm_reduce_ms33 & multm_reduce_mc32;
  assign multm_reduce_add3b1_maj3b_xy23 = multm_reduce_ms34 & multm_reduce_mc33;
  assign multm_reduce_add3b1_maj3b_xy24 = multm_reduce_ms35 & multm_reduce_mc34;
  assign multm_reduce_add3b1_maj3b_xy25 = multm_reduce_ms36 & multm_reduce_mc35;
  assign multm_reduce_add3b1_maj3b_xy26 = multm_reduce_ms37 & multm_reduce_mc36;
  assign multm_reduce_add3b1_maj3b_xy27 = multm_reduce_ms38 & multm_reduce_mc37;
  assign multm_reduce_add3b1_maj3b_xy28 = multm_reduce_ms39 & multm_reduce_mc38;
  assign multm_reduce_add3b1_maj3b_xy29 = multm_reduce_ms40 & multm_reduce_mc39;
  assign multm_reduce_add3b1_maj3b_xy30 = multm_reduce_ms41 & multm_reduce_mc40;
  assign multm_reduce_add3b1_maj3b_xy31 = multm_reduce_ms42 & multm_reduce_mc41;
  assign multm_reduce_add3b1_maj3b_xy32 = multm_reduce_ms43 & multm_reduce_mc42;
  assign multm_reduce_add3b1_maj3b_xy33 = multm_reduce_ms44 & multm_reduce_mc43;
  assign multm_reduce_add3b1_maj3b_xy34 = multm_reduce_ms45 & multm_reduce_mc44;
  assign multm_reduce_add3b1_maj3b_xy35 = multm_reduce_ms46 & multm_reduce_mc45;
  assign multm_reduce_add3b1_maj3b_xy36 = multm_reduce_ms47 & multm_reduce_mc46;
  assign multm_reduce_add3b1_maj3b_xy37 = multm_reduce_ms48 & multm_reduce_mc47;
  assign multm_reduce_add3b1_maj3b_xy38 = multm_reduce_ms49 & multm_reduce_mc48;
  assign multm_reduce_add3b1_maj3b_xy39 = multm_reduce_ms50 & multm_reduce_mc49;
  assign multm_reduce_add3b1_maj3b_xy40 = multm_reduce_ms51 & multm_reduce_mc50;
  assign multm_reduce_add3b1_maj3b_xy41 = multm_reduce_ms52 & multm_reduce_mc51;
  assign multm_reduce_add3b1_maj3b_xy42 = multm_reduce_ms53 & multm_reduce_mc52;
  assign multm_reduce_add3b1_maj3b_xy43 = multm_reduce_ms54 & multm_reduce_mc53;
  assign multm_reduce_add3b1_maj3b_xy44 = multm_reduce_ms55 & multm_reduce_mc54;
  assign multm_reduce_add3b1_maj3b_xy45 = multm_reduce_ms56 & multm_reduce_mc55;
  assign multm_reduce_add3b1_maj3b_xy46 = multm_reduce_ms57 & multm_reduce_mc56;
  assign multm_reduce_add3b1_maj3b_xy47 = multm_reduce_ms58 & multm_reduce_mc57;
  assign multm_reduce_add3b1_maj3b_xy48 = multm_reduce_ms59 & multm_reduce_mc58;
  assign multm_reduce_add3b1_maj3b_xy49 = multm_reduce_ms60 & multm_reduce_mc59;
  assign multm_reduce_add3b1_maj3b_xy50 = multm_reduce_ms61 & multm_reduce_mc60;
  assign multm_reduce_add3b1_maj3b_xy51 = multm_reduce_ms62 & multm_reduce_mc61;
  assign multm_reduce_add3b1_maj3b_xy52 = multm_reduce_ms63 & multm_reduce_mc62;
  assign multm_reduce_add3b1_maj3b_xy53 = multm_reduce_ms64 & multm_reduce_mc63;
  assign multm_reduce_add3b1_maj3b_xy54 = multm_reduce_ms65 & multm_reduce_mc64;
  assign multm_reduce_add3b1_maj3b_xy55 = multm_reduce_ms66 & multm_reduce_mc65;
  assign multm_reduce_add3b1_maj3b_xy56 = multm_reduce_ms67 & multm_reduce_mc66;
  assign multm_reduce_add3b1_maj3b_xy57 = multm_reduce_ms68 & multm_reduce_mc67;
  assign multm_reduce_add3b1_maj3b_xy58 = multm_reduce_ms69 & multm_reduce_mc68;
  assign multm_reduce_add3b1_maj3b_xy59 = multm_reduce_ms70 & multm_reduce_mc69;
  assign multm_reduce_add3b1_maj3b_xy60 = multm_reduce_ms71 & multm_reduce_mc70;
  assign multm_reduce_add3b1_maj3b_xy61 = multm_reduce_ms72 & multm_reduce_mc71;
  assign multm_reduce_add3b1_maj3b_xy62 = multm_reduce_ms73 & multm_reduce_mc72;
  assign multm_reduce_add3b1_maj3b_xy63 = multm_reduce_ms74 & multm_reduce_mc73;
  assign multm_reduce_add3b1_maj3b_xy64 = multm_reduce_ms75 & multm_reduce_mc74;
  assign multm_reduce_add3b1_maj3b_xy65 = multm_reduce_ms76 & multm_reduce_mc75;
  assign multm_reduce_add3b1_maj3b_xy66 = multm_reduce_ms77 & multm_reduce_mc76;
  assign multm_reduce_add3b1_maj3b_xy67 = multm_reduce_ms78 & multm_reduce_mc77;
  assign multm_reduce_add3b1_maj3b_xy68 = multm_reduce_ms79 & multm_reduce_mc78;
  assign multm_reduce_add3b1_maj3b_xy69 = multm_reduce_ms80 & multm_reduce_mc79;
  assign multm_reduce_add3b1_maj3b_xy70 = multm_reduce_ms81 & multm_reduce_mc80;
  assign multm_reduce_add3b1_maj3b_xy71 = multm_reduce_ms82 & multm_reduce_mc81;
  assign multm_reduce_add3b1_maj3b_xy72 = multm_reduce_ms83 & multm_reduce_mc82;
  assign multm_reduce_add3b1_maj3b_xy73 = multm_reduce_ms84 & multm_reduce_mc83;
  assign multm_reduce_add3b1_maj3b_xy74 = multm_reduce_ms85 & multm_reduce_mc84;
  assign multm_reduce_add3b1_maj3b_xy75 = multm_reduce_ms86 & multm_reduce_mc85;
  assign multm_reduce_add3b1_maj3b_xy76 = multm_reduce_ms87 & multm_reduce_mc86;
  assign multm_reduce_add3b1_maj3b_xy77 = multm_reduce_ms88 & multm_reduce_mc87;
  assign multm_reduce_add3b1_maj3b_xy78 = multm_reduce_ms89 & multm_reduce_mc88;
  assign multm_reduce_add3b1_maj3b_xy79 = multm_reduce_ms90 & multm_reduce_mc89;
  assign multm_reduce_add3b1_maj3b_xy80 = multm_reduce_ms91 & multm_reduce_mc90;
  assign multm_reduce_add3b1_maj3b_xy81 = multm_reduce_ms92 & multm_reduce_mc91;
  assign multm_reduce_add3b1_maj3b_xy82 = multm_reduce_ms93 & multm_reduce_mc92;
  assign multm_reduce_add3b1_maj3b_xy83 = multm_reduce_ms94 & multm_reduce_mc93;
  assign multm_reduce_add3b1_maj3b_xy84 = multm_reduce_ms95 & multm_reduce_mc94;
  assign multm_reduce_add3b1_maj3b_xy85 = multm_reduce_ms96 & multm_reduce_mc95;
  assign multm_reduce_add3b1_maj3b_xy86 = multm_reduce_ms97 & multm_reduce_mc96;
  assign multm_reduce_add3b1_maj3b_xy87 = multm_reduce_ms98 & multm_reduce_mc97;
  assign multm_reduce_add3b1_maj3b_xy88 = multm_reduce_ms99 & multm_reduce_mc98;
  assign multm_reduce_add3b1_maj3b_xy89 = multm_reduce_ms100 & multm_reduce_mc99;
  assign multm_reduce_add3b1_maj3b_xy90 = multm_reduce_ms101 & multm_reduce_mc100;
  assign multm_reduce_add3b1_maj3b_xy91 = multm_reduce_ms102 & multm_reduce_mc101;
  assign multm_reduce_add3b1_maj3b_xy92 = multm_reduce_ms103 & multm_reduce_mc102;
  assign multm_reduce_add3b1_maj3b_xy93 = multm_reduce_ms104 & multm_reduce_mc103;
  assign multm_reduce_add3b1_maj3b_xy94 = multm_reduce_ms105 & multm_reduce_mc104;
  assign multm_reduce_add3b1_maj3b_xy95 = multm_reduce_ms106 & multm_reduce_mc105;
  assign multm_reduce_add3b1_maj3b_xy96 = multm_reduce_ms107 & multm_reduce_mc106;
  assign multm_reduce_add3b1_maj3b_xy97 = multm_reduce_ms108 & multm_reduce_mc107;
  assign multm_reduce_add3b1_maj3b_xy98 = multm_reduce_ms109 & multm_reduce_mc108;
  assign multm_reduce_add3b1_maj3b_xy99 = multm_reduce_ms110 & multm_reduce_mc109;
  assign multm_reduce_add3b1_maj3b_xy100 = multm_reduce_ms111 & multm_reduce_mc110;
  assign multm_reduce_add3b1_maj3b_xy101 = multm_reduce_ms112 & multm_reduce_mc111;
  assign multm_reduce_add3b1_maj3b_xy102 = multm_reduce_ms113 & multm_reduce_mc112;
  assign multm_reduce_add3b1_maj3b_xy103 = multm_reduce_ms114 & multm_reduce_mc113;
  assign multm_reduce_add3b1_maj3b_xy104 = multm_reduce_ms115 & multm_reduce_mc114;
  assign multm_reduce_add3b1_maj3b_xy105 = multm_reduce_ms116 & multm_reduce_mc115;
  assign multm_reduce_add3b1_maj3b_xy106 = multm_reduce_ms117 & multm_reduce_mc116;
  assign multm_reduce_add3b1_maj3b_xy107 = multm_reduce_ms118 & multm_reduce_mc117;
  assign multm_reduce_add3b1_maj3b_xy108 = multm_reduce_ms119 & multm_reduce_mc118;
  assign multm_reduce_add3b1_maj3b_xy109 = multm_reduce_ms120 & multm_reduce_mc119;
  assign multm_reduce_add3b1_maj3b_xy110 = multm_reduce_ms121 & multm_reduce_mc120;
  assign multm_reduce_add3b1_maj3b_xy111 = multm_reduce_ms122 & multm_reduce_mc121;
  assign multm_reduce_add3b1_maj3b_xy112 = multm_reduce_ms123 & multm_reduce_mc122;
  assign multm_reduce_add3b1_maj3b_xy113 = multm_reduce_ms124 & multm_reduce_mc123;
  assign multm_reduce_add3b1_maj3b_xy114 = multm_reduce_ms125 & multm_reduce_mc124;
  assign multm_reduce_add3b1_maj3b_xy115 = multm_reduce_ms126 & multm_reduce_mc125;
  assign multm_reduce_add3b1_maj3b_xy116 = multm_reduce_ms127 & multm_reduce_mc126;
  assign multm_reduce_add3b1_maj3b_xy117 = multm_reduce_ms128 & multm_reduce_mc127;
  assign multm_reduce_add3b1_maj3b_xy118 = multm_reduce_ms129 & multm_reduce_mc128;
  assign multm_reduce_add3b1_maj3b_xy119 = multm_reduce_ms130 & multm_reduce_mc129;
  assign multm_reduce_add3b1_maj3b_xy120 = multm_reduce_ms131 & multm_reduce_mc130;
  assign multm_reduce_add3b1_maj3b_xy121 = multm_reduce_ms132 & multm_reduce_mc131;
  assign multm_reduce_add3b1_maj3b_xy122 = multm_reduce_ms133 & multm_reduce_mc132;
  assign multm_reduce_add3b1_maj3b_xy123 = multm_reduce_ms134 & multm_reduce_mc133;
  assign multm_reduce_add3b1_maj3b_xy124 = multm_reduce_ms135 & multm_reduce_mc134;
  assign multm_reduce_add3b1_maj3b_xy125 = multm_reduce_ms136 & multm_reduce_mc135;
  assign multm_reduce_add3b1_maj3b_xy126 = multm_reduce_ms137 & multm_reduce_mc136;
  assign multm_reduce_add3b1_maj3b_xy127 = multm_reduce_ms138 & multm_reduce_mc137;
  assign multm_reduce_add3b1_maj3b_xy128 = multm_reduce_ms139 & multm_reduce_mc138;
  assign multm_reduce_add3b1_maj3b_xy129 = multm_reduce_ms140 & multm_reduce_mc139;
  assign multm_reduce_add3b1_maj3b_xy130 = multm_reduce_ms141 & multm_reduce_mc140;
  assign multm_reduce_add3b1_maj3b_xy131 = multm_reduce_ms142 & multm_reduce_mc141;
  assign multm_reduce_add3b1_maj3b_xy132 = multm_reduce_ms143 & multm_reduce_mc142;
  assign multm_reduce_add3b1_maj3b_xy133 = multm_reduce_ms144 & multm_reduce_mc143;
  assign multm_reduce_add3b1_maj3b_xy134 = multm_reduce_ms145 & multm_reduce_mc144;
  assign multm_reduce_add3b1_maj3b_xy135 = multm_reduce_ms146 & multm_reduce_mc145;
  assign multm_reduce_add3b1_maj3b_xy136 = multm_reduce_ms147 & multm_reduce_mc146;
  assign multm_reduce_add3b1_maj3b_xy137 = multm_reduce_ms148 & multm_reduce_mc147;
  assign multm_reduce_add3b1_maj3b_xy138 = multm_reduce_ms149 & multm_reduce_mc148;
  assign multm_reduce_add3b1_maj3b_xy139 = multm_reduce_ms150 & multm_reduce_mc149;
  assign multm_reduce_add3b1_maj3b_xy140 = multm_reduce_ms151 & multm_reduce_mc150;
  assign multm_reduce_add3b1_maj3b_xy141 = multm_reduce_ms152 & multm_reduce_mc151;
  assign multm_reduce_add3b1_maj3b_xy142 = multm_reduce_ms153 & multm_reduce_mc152;
  assign multm_reduce_add3b1_maj3b_xy143 = multm_reduce_ms154 & multm_reduce_mc153;
  assign multm_reduce_add3b1_maj3b_xy144 = multm_reduce_ms155 & multm_reduce_mc154;
  assign multm_reduce_add3b1_maj3b_xy145 = multm_reduce_ms156 & multm_reduce_mc155;
  assign multm_reduce_add3b1_maj3b_xy146 = multm_reduce_ms157 & multm_reduce_mc156;
  assign multm_reduce_add3b1_maj3b_xy147 = multm_reduce_ms158 & multm_reduce_mc157;
  assign multm_reduce_add3b1_maj3b_xy148 = multm_reduce_ms159 & multm_reduce_mc158;
  assign multm_reduce_add3b1_maj3b_xy149 = multm_reduce_ms160 & multm_reduce_mc159;
  assign multm_reduce_add3b1_maj3b_xy150 = multm_reduce_ms161 & multm_reduce_mc160;
  assign multm_reduce_add3b1_maj3b_xy151 = multm_reduce_ms162 & multm_reduce_mc161;
  assign multm_reduce_add3b1_maj3b_xy152 = multm_reduce_ms163 & multm_reduce_mc162;
  assign multm_reduce_add3b1_maj3b_xy153 = multm_reduce_ms164 & multm_reduce_mc163;
  assign multm_reduce_add3b1_maj3b_xy154 = multm_reduce_ms165 & multm_reduce_mc164;
  assign multm_reduce_add3b1_maj3b_xy155 = multm_reduce_ms166 & multm_reduce_mc165;
  assign multm_reduce_add3b1_maj3b_xy156 = multm_reduce_ms167 & multm_reduce_mc166;
  assign multm_reduce_add3b1_maj3b_xy157 = multm_reduce_ms168 & multm_reduce_mc167;
  assign multm_reduce_add3b1_maj3b_xy158 = multm_reduce_ms169 & multm_reduce_mc168;
  assign multm_reduce_add3b1_maj3b_xy159 = multm_reduce_ms170 & multm_reduce_mc169;
  assign multm_reduce_add3b1_maj3b_xy160 = multm_reduce_ms171 & multm_reduce_mc170;
  assign multm_reduce_add3b1_maj3b_xy161 = multm_reduce_ms172 & multm_reduce_mc171;
  assign multm_reduce_add3b1_maj3b_xy162 = multm_reduce_ms173 & multm_reduce_mc172;
  assign multm_reduce_add3b1_maj3b_xy163 = multm_reduce_ms174 & multm_reduce_mc173;
  assign multm_reduce_add3b1_maj3b_xy164 = multm_reduce_ms175 & multm_reduce_mc174;
  assign multm_reduce_add3b1_maj3b_xy165 = multm_reduce_ms176 & multm_reduce_mc175;
  assign multm_reduce_add3b1_maj3b_xy166 = multm_reduce_ms177 & multm_reduce_mc176;
  assign multm_reduce_add3b1_maj3b_xy167 = multm_reduce_ms178 & multm_reduce_mc177;
  assign multm_reduce_add3b1_maj3b_xy168 = multm_reduce_ms179 & multm_reduce_mc178;
  assign multm_reduce_add3b1_maj3b_xy169 = multm_reduce_ms180 & multm_reduce_mc179;
  assign multm_reduce_add3b1_maj3b_xy170 = multm_reduce_ms181 & multm_reduce_mc180;
  assign multm_reduce_add3b1_maj3b_xy171 = multm_reduce_ms182 & multm_reduce_mc181;
  assign multm_reduce_add3b1_maj3b_xy172 = multm_reduce_ms183 & multm_reduce_mc182;
  assign multm_reduce_add3b1_xor3b_wx0 = multm_reduce_sb0 ^ multm_reduce_ms11;
  assign multm_reduce_add3b1_xor3b_wx1 = multm_reduce_sb1 ^ multm_reduce_ms12;
  assign multm_reduce_add3b1_xor3b_wx2 = multm_reduce_sb2 ^ multm_reduce_ms13;
  assign multm_reduce_add3b1_xor3b_wx3 = multm_reduce_sb3 ^ multm_reduce_ms14;
  assign multm_reduce_add3b1_xor3b_wx4 = multm_reduce_sb4 ^ multm_reduce_ms15;
  assign multm_reduce_add3b1_xor3b_wx5 = multm_reduce_sb5 ^ multm_reduce_ms16;
  assign multm_reduce_add3b1_xor3b_wx6 = multm_reduce_sb6 ^ multm_reduce_ms17;
  assign multm_reduce_add3b1_xor3b_wx7 = multm_reduce_sb7 ^ multm_reduce_ms18;
  assign multm_reduce_add3b1_xor3b_wx8 = multm_reduce_sb8 ^ multm_reduce_ms19;
  assign multm_reduce_add3b1_xor3b_wx9 = multm_reduce_sb9 ^ multm_reduce_ms20;
  assign multm_reduce_add3b1_xor3b_wx10 = multm_reduce_sb10 ^ multm_reduce_ms21;
  assign multm_reduce_add3b1_xor3b_wx11 = multm_reduce_sb11 ^ multm_reduce_ms22;
  assign multm_reduce_add3b1_xor3b_wx12 = multm_reduce_sb12 ^ multm_reduce_ms23;
  assign multm_reduce_add3b1_xor3b_wx13 = multm_reduce_sb13 ^ multm_reduce_ms24;
  assign multm_reduce_add3b1_xor3b_wx14 = multm_reduce_sb14 ^ multm_reduce_ms25;
  assign multm_reduce_add3b1_xor3b_wx15 = multm_reduce_sb15 ^ multm_reduce_ms26;
  assign multm_reduce_add3b1_xor3b_wx16 = multm_reduce_sb16 ^ multm_reduce_ms27;
  assign multm_reduce_add3b1_xor3b_wx17 = multm_reduce_sb17 ^ multm_reduce_ms28;
  assign multm_reduce_add3b1_xor3b_wx18 = multm_reduce_sb18 ^ multm_reduce_ms29;
  assign multm_reduce_add3b1_xor3b_wx19 = multm_reduce_sb19 ^ multm_reduce_ms30;
  assign multm_reduce_add3b1_xor3b_wx20 = multm_reduce_sb20 ^ multm_reduce_ms31;
  assign multm_reduce_add3b1_xor3b_wx21 = multm_reduce_sb21 ^ multm_reduce_ms32;
  assign multm_reduce_add3b1_xor3b_wx22 = multm_reduce_sb22 ^ multm_reduce_ms33;
  assign multm_reduce_add3b1_xor3b_wx23 = multm_reduce_sb23 ^ multm_reduce_ms34;
  assign multm_reduce_add3b1_xor3b_wx24 = multm_reduce_sb24 ^ multm_reduce_ms35;
  assign multm_reduce_add3b1_xor3b_wx25 = multm_reduce_sb25 ^ multm_reduce_ms36;
  assign multm_reduce_add3b1_xor3b_wx26 = multm_reduce_sb26 ^ multm_reduce_ms37;
  assign multm_reduce_add3b1_xor3b_wx27 = multm_reduce_sb27 ^ multm_reduce_ms38;
  assign multm_reduce_add3b1_xor3b_wx28 = multm_reduce_sb28 ^ multm_reduce_ms39;
  assign multm_reduce_add3b1_xor3b_wx29 = multm_reduce_sb29 ^ multm_reduce_ms40;
  assign multm_reduce_add3b1_xor3b_wx30 = multm_reduce_sb30 ^ multm_reduce_ms41;
  assign multm_reduce_add3b1_xor3b_wx31 = multm_reduce_sb31 ^ multm_reduce_ms42;
  assign multm_reduce_add3b1_xor3b_wx32 = multm_reduce_sb32 ^ multm_reduce_ms43;
  assign multm_reduce_add3b1_xor3b_wx33 = multm_reduce_sb33 ^ multm_reduce_ms44;
  assign multm_reduce_add3b1_xor3b_wx34 = multm_reduce_sb34 ^ multm_reduce_ms45;
  assign multm_reduce_add3b1_xor3b_wx35 = multm_reduce_sb35 ^ multm_reduce_ms46;
  assign multm_reduce_add3b1_xor3b_wx36 = multm_reduce_sb36 ^ multm_reduce_ms47;
  assign multm_reduce_add3b1_xor3b_wx37 = multm_reduce_sb37 ^ multm_reduce_ms48;
  assign multm_reduce_add3b1_xor3b_wx38 = multm_reduce_sb38 ^ multm_reduce_ms49;
  assign multm_reduce_add3b1_xor3b_wx39 = multm_reduce_sb39 ^ multm_reduce_ms50;
  assign multm_reduce_add3b1_xor3b_wx40 = multm_reduce_sb40 ^ multm_reduce_ms51;
  assign multm_reduce_add3b1_xor3b_wx41 = multm_reduce_sb41 ^ multm_reduce_ms52;
  assign multm_reduce_add3b1_xor3b_wx42 = multm_reduce_sb42 ^ multm_reduce_ms53;
  assign multm_reduce_add3b1_xor3b_wx43 = multm_reduce_sb43 ^ multm_reduce_ms54;
  assign multm_reduce_add3b1_xor3b_wx44 = multm_reduce_sb44 ^ multm_reduce_ms55;
  assign multm_reduce_add3b1_xor3b_wx45 = multm_reduce_sb45 ^ multm_reduce_ms56;
  assign multm_reduce_add3b1_xor3b_wx46 = multm_reduce_sb46 ^ multm_reduce_ms57;
  assign multm_reduce_add3b1_xor3b_wx47 = multm_reduce_sb47 ^ multm_reduce_ms58;
  assign multm_reduce_add3b1_xor3b_wx48 = multm_reduce_sb48 ^ multm_reduce_ms59;
  assign multm_reduce_add3b1_xor3b_wx49 = multm_reduce_sb49 ^ multm_reduce_ms60;
  assign multm_reduce_add3b1_xor3b_wx50 = multm_reduce_sb50 ^ multm_reduce_ms61;
  assign multm_reduce_add3b1_xor3b_wx51 = multm_reduce_sb51 ^ multm_reduce_ms62;
  assign multm_reduce_add3b1_xor3b_wx52 = multm_reduce_sb52 ^ multm_reduce_ms63;
  assign multm_reduce_add3b1_xor3b_wx53 = multm_reduce_sb53 ^ multm_reduce_ms64;
  assign multm_reduce_add3b1_xor3b_wx54 = multm_reduce_sb54 ^ multm_reduce_ms65;
  assign multm_reduce_add3b1_xor3b_wx55 = multm_reduce_sb55 ^ multm_reduce_ms66;
  assign multm_reduce_add3b1_xor3b_wx56 = multm_reduce_sb56 ^ multm_reduce_ms67;
  assign multm_reduce_add3b1_xor3b_wx57 = multm_reduce_sb57 ^ multm_reduce_ms68;
  assign multm_reduce_add3b1_xor3b_wx58 = multm_reduce_sb58 ^ multm_reduce_ms69;
  assign multm_reduce_add3b1_xor3b_wx59 = multm_reduce_sb59 ^ multm_reduce_ms70;
  assign multm_reduce_add3b1_xor3b_wx60 = multm_reduce_sb60 ^ multm_reduce_ms71;
  assign multm_reduce_add3b1_xor3b_wx61 = multm_reduce_sb61 ^ multm_reduce_ms72;
  assign multm_reduce_add3b1_xor3b_wx62 = multm_reduce_sb62 ^ multm_reduce_ms73;
  assign multm_reduce_add3b1_xor3b_wx63 = multm_reduce_sb63 ^ multm_reduce_ms74;
  assign multm_reduce_add3b1_xor3b_wx64 = multm_reduce_sb64 ^ multm_reduce_ms75;
  assign multm_reduce_add3b1_xor3b_wx65 = multm_reduce_sb65 ^ multm_reduce_ms76;
  assign multm_reduce_add3b1_xor3b_wx66 = multm_reduce_sb66 ^ multm_reduce_ms77;
  assign multm_reduce_add3b1_xor3b_wx67 = multm_reduce_sb67 ^ multm_reduce_ms78;
  assign multm_reduce_add3b1_xor3b_wx68 = multm_reduce_sb68 ^ multm_reduce_ms79;
  assign multm_reduce_add3b1_xor3b_wx69 = multm_reduce_sb69 ^ multm_reduce_ms80;
  assign multm_reduce_add3b1_xor3b_wx70 = multm_reduce_sb70 ^ multm_reduce_ms81;
  assign multm_reduce_add3b1_xor3b_wx71 = multm_reduce_sb71 ^ multm_reduce_ms82;
  assign multm_reduce_add3b1_xor3b_wx72 = multm_reduce_sb72 ^ multm_reduce_ms83;
  assign multm_reduce_add3b1_xor3b_wx73 = multm_reduce_sb73 ^ multm_reduce_ms84;
  assign multm_reduce_add3b1_xor3b_wx74 = multm_reduce_sb74 ^ multm_reduce_ms85;
  assign multm_reduce_add3b1_xor3b_wx75 = multm_reduce_sb75 ^ multm_reduce_ms86;
  assign multm_reduce_add3b1_xor3b_wx76 = multm_reduce_sb76 ^ multm_reduce_ms87;
  assign multm_reduce_add3b1_xor3b_wx77 = multm_reduce_sb77 ^ multm_reduce_ms88;
  assign multm_reduce_add3b1_xor3b_wx78 = multm_reduce_sb78 ^ multm_reduce_ms89;
  assign multm_reduce_add3b1_xor3b_wx79 = multm_reduce_sb79 ^ multm_reduce_ms90;
  assign multm_reduce_add3b1_xor3b_wx80 = multm_reduce_sb80 ^ multm_reduce_ms91;
  assign multm_reduce_add3b1_xor3b_wx81 = multm_reduce_sb81 ^ multm_reduce_ms92;
  assign multm_reduce_add3b1_xor3b_wx82 = multm_reduce_sb82 ^ multm_reduce_ms93;
  assign multm_reduce_add3b1_xor3b_wx83 = multm_reduce_sb83 ^ multm_reduce_ms94;
  assign multm_reduce_add3b1_xor3b_wx84 = multm_reduce_sb84 ^ multm_reduce_ms95;
  assign multm_reduce_add3b1_xor3b_wx85 = multm_reduce_sb85 ^ multm_reduce_ms96;
  assign multm_reduce_add3b1_xor3b_wx86 = multm_reduce_sb86 ^ multm_reduce_ms97;
  assign multm_reduce_add3b1_xor3b_wx87 = multm_reduce_sb87 ^ multm_reduce_ms98;
  assign multm_reduce_add3b1_xor3b_wx88 = multm_reduce_sb88 ^ multm_reduce_ms99;
  assign multm_reduce_add3b1_xor3b_wx89 = multm_reduce_sb89 ^ multm_reduce_ms100;
  assign multm_reduce_add3b1_xor3b_wx90 = multm_reduce_sb90 ^ multm_reduce_ms101;
  assign multm_reduce_add3b1_xor3b_wx91 = multm_reduce_sb91 ^ multm_reduce_ms102;
  assign multm_reduce_add3b1_xor3b_wx92 = multm_reduce_sb92 ^ multm_reduce_ms103;
  assign multm_reduce_add3b1_xor3b_wx93 = multm_reduce_sb93 ^ multm_reduce_ms104;
  assign multm_reduce_add3b1_xor3b_wx94 = multm_reduce_sb94 ^ multm_reduce_ms105;
  assign multm_reduce_add3b1_xor3b_wx95 = multm_reduce_sb95 ^ multm_reduce_ms106;
  assign multm_reduce_add3b1_xor3b_wx96 = multm_reduce_sb96 ^ multm_reduce_ms107;
  assign multm_reduce_add3b1_xor3b_wx97 = multm_reduce_sb97 ^ multm_reduce_ms108;
  assign multm_reduce_add3b1_xor3b_wx98 = multm_reduce_sb98 ^ multm_reduce_ms109;
  assign multm_reduce_add3b1_xor3b_wx99 = multm_reduce_sb99 ^ multm_reduce_ms110;
  assign multm_reduce_add3b1_xor3b_wx100 = multm_reduce_sb100 ^ multm_reduce_ms111;
  assign multm_reduce_add3b1_xor3b_wx101 = multm_reduce_sb101 ^ multm_reduce_ms112;
  assign multm_reduce_add3b1_xor3b_wx102 = multm_reduce_sb102 ^ multm_reduce_ms113;
  assign multm_reduce_add3b1_xor3b_wx103 = multm_reduce_sb103 ^ multm_reduce_ms114;
  assign multm_reduce_add3b1_xor3b_wx104 = multm_reduce_sb104 ^ multm_reduce_ms115;
  assign multm_reduce_add3b1_xor3b_wx105 = multm_reduce_sb105 ^ multm_reduce_ms116;
  assign multm_reduce_add3b1_xor3b_wx106 = multm_reduce_sb106 ^ multm_reduce_ms117;
  assign multm_reduce_add3b1_xor3b_wx107 = multm_reduce_sb107 ^ multm_reduce_ms118;
  assign multm_reduce_add3b1_xor3b_wx108 = multm_reduce_sb108 ^ multm_reduce_ms119;
  assign multm_reduce_add3b1_xor3b_wx109 = multm_reduce_sb109 ^ multm_reduce_ms120;
  assign multm_reduce_add3b1_xor3b_wx110 = multm_reduce_sb110 ^ multm_reduce_ms121;
  assign multm_reduce_add3b1_xor3b_wx111 = multm_reduce_sb111 ^ multm_reduce_ms122;
  assign multm_reduce_add3b1_xor3b_wx112 = multm_reduce_sb112 ^ multm_reduce_ms123;
  assign multm_reduce_add3b1_xor3b_wx113 = multm_reduce_sb113 ^ multm_reduce_ms124;
  assign multm_reduce_add3b1_xor3b_wx114 = multm_reduce_sb114 ^ multm_reduce_ms125;
  assign multm_reduce_add3b1_xor3b_wx115 = multm_reduce_sb115 ^ multm_reduce_ms126;
  assign multm_reduce_add3b1_xor3b_wx116 = multm_reduce_sb116 ^ multm_reduce_ms127;
  assign multm_reduce_add3b1_xor3b_wx117 = multm_reduce_sb117 ^ multm_reduce_ms128;
  assign multm_reduce_add3b1_xor3b_wx118 = multm_reduce_sb118 ^ multm_reduce_ms129;
  assign multm_reduce_add3b1_xor3b_wx119 = multm_reduce_sb119 ^ multm_reduce_ms130;
  assign multm_reduce_add3b1_xor3b_wx120 = multm_reduce_sb120 ^ multm_reduce_ms131;
  assign multm_reduce_add3b1_xor3b_wx121 = multm_reduce_sb121 ^ multm_reduce_ms132;
  assign multm_reduce_add3b1_xor3b_wx122 = multm_reduce_sb122 ^ multm_reduce_ms133;
  assign multm_reduce_add3b1_xor3b_wx123 = multm_reduce_sb123 ^ multm_reduce_ms134;
  assign multm_reduce_add3b1_xor3b_wx124 = multm_reduce_sb124 ^ multm_reduce_ms135;
  assign multm_reduce_add3b1_xor3b_wx125 = multm_reduce_sb125 ^ multm_reduce_ms136;
  assign multm_reduce_add3b1_xor3b_wx126 = multm_reduce_sb126 ^ multm_reduce_ms137;
  assign multm_reduce_add3b1_xor3b_wx127 = multm_reduce_sb127 ^ multm_reduce_ms138;
  assign multm_reduce_add3b1_xor3b_wx128 = multm_reduce_sb128 ^ multm_reduce_ms139;
  assign multm_reduce_add3b1_xor3b_wx129 = multm_reduce_sb129 ^ multm_reduce_ms140;
  assign multm_reduce_add3b1_xor3b_wx130 = multm_reduce_sb130 ^ multm_reduce_ms141;
  assign multm_reduce_add3b1_xor3b_wx131 = multm_reduce_sb131 ^ multm_reduce_ms142;
  assign multm_reduce_add3b1_xor3b_wx132 = multm_reduce_sb132 ^ multm_reduce_ms143;
  assign multm_reduce_add3b1_xor3b_wx133 = multm_reduce_sb133 ^ multm_reduce_ms144;
  assign multm_reduce_add3b1_xor3b_wx134 = multm_reduce_sb134 ^ multm_reduce_ms145;
  assign multm_reduce_add3b1_xor3b_wx135 = multm_reduce_sb135 ^ multm_reduce_ms146;
  assign multm_reduce_add3b1_xor3b_wx136 = multm_reduce_sb136 ^ multm_reduce_ms147;
  assign multm_reduce_add3b1_xor3b_wx137 = multm_reduce_sb137 ^ multm_reduce_ms148;
  assign multm_reduce_add3b1_xor3b_wx138 = multm_reduce_sb138 ^ multm_reduce_ms149;
  assign multm_reduce_add3b1_xor3b_wx139 = multm_reduce_sb139 ^ multm_reduce_ms150;
  assign multm_reduce_add3b1_xor3b_wx140 = multm_reduce_sb140 ^ multm_reduce_ms151;
  assign multm_reduce_add3b1_xor3b_wx141 = multm_reduce_sb141 ^ multm_reduce_ms152;
  assign multm_reduce_add3b1_xor3b_wx142 = multm_reduce_sb142 ^ multm_reduce_ms153;
  assign multm_reduce_add3b1_xor3b_wx143 = multm_reduce_sb143 ^ multm_reduce_ms154;
  assign multm_reduce_add3b1_xor3b_wx144 = multm_reduce_sb144 ^ multm_reduce_ms155;
  assign multm_reduce_add3b1_xor3b_wx145 = multm_reduce_sb145 ^ multm_reduce_ms156;
  assign multm_reduce_add3b1_xor3b_wx146 = multm_reduce_sb146 ^ multm_reduce_ms157;
  assign multm_reduce_add3b1_xor3b_wx147 = multm_reduce_sb147 ^ multm_reduce_ms158;
  assign multm_reduce_add3b1_xor3b_wx148 = multm_reduce_sb148 ^ multm_reduce_ms159;
  assign multm_reduce_add3b1_xor3b_wx149 = multm_reduce_sb149 ^ multm_reduce_ms160;
  assign multm_reduce_add3b1_xor3b_wx150 = multm_reduce_sb150 ^ multm_reduce_ms161;
  assign multm_reduce_add3b1_xor3b_wx151 = multm_reduce_sb151 ^ multm_reduce_ms162;
  assign multm_reduce_add3b1_xor3b_wx152 = multm_reduce_sb152 ^ multm_reduce_ms163;
  assign multm_reduce_add3b1_xor3b_wx153 = multm_reduce_sb153 ^ multm_reduce_ms164;
  assign multm_reduce_add3b1_xor3b_wx154 = multm_reduce_sb154 ^ multm_reduce_ms165;
  assign multm_reduce_add3b1_xor3b_wx155 = multm_reduce_sb155 ^ multm_reduce_ms166;
  assign multm_reduce_add3b1_xor3b_wx156 = multm_reduce_sb156 ^ multm_reduce_ms167;
  assign multm_reduce_add3b1_xor3b_wx157 = multm_reduce_sb157 ^ multm_reduce_ms168;
  assign multm_reduce_add3b1_xor3b_wx158 = multm_reduce_sb158 ^ multm_reduce_ms169;
  assign multm_reduce_add3b1_xor3b_wx159 = multm_reduce_sb159 ^ multm_reduce_ms170;
  assign multm_reduce_add3b1_xor3b_wx160 = multm_reduce_sb160 ^ multm_reduce_ms171;
  assign multm_reduce_add3b1_xor3b_wx161 = multm_reduce_sb161 ^ multm_reduce_ms172;
  assign multm_reduce_add3b1_xor3b_wx162 = multm_reduce_sb162 ^ multm_reduce_ms173;
  assign multm_reduce_add3b1_xor3b_wx163 = multm_reduce_sb163 ^ multm_reduce_ms174;
  assign multm_reduce_add3b1_xor3b_wx164 = multm_reduce_sb164 ^ multm_reduce_ms175;
  assign multm_reduce_add3b1_xor3b_wx165 = multm_reduce_sb165 ^ multm_reduce_ms176;
  assign multm_reduce_add3b1_xor3b_wx166 = multm_reduce_sb166 ^ multm_reduce_ms177;
  assign multm_reduce_add3b1_xor3b_wx167 = multm_reduce_sb167 ^ multm_reduce_ms178;
  assign multm_reduce_add3b1_xor3b_wx168 = multm_reduce_sb168 ^ multm_reduce_ms179;
  assign multm_reduce_add3b1_xor3b_wx169 = multm_reduce_sb169 ^ multm_reduce_ms180;
  assign multm_reduce_add3b1_xor3b_wx170 = multm_reduce_sb170 ^ multm_reduce_ms181;
  assign multm_reduce_add3b1_xor3b_wx171 = multm_reduce_sb171 ^ multm_reduce_ms182;
  assign multm_reduce_add3b1_xor3b_wx172 = multm_reduce_sb172 ^ multm_reduce_ms183;
  assign multm_reduce_mc10 = multm_reduce_add3b0_maj3b_or3b_wx10 | multm_reduce_add3b0_maj3b_xy10;
  assign multm_reduce_mc11 = multm_reduce_add3b0_maj3b_or3b_wx11 | multm_reduce_add3b0_maj3b_xy11;
  assign multm_reduce_mc12 = multm_reduce_add3b0_maj3b_or3b_wx12 | multm_reduce_add3b0_maj3b_xy12;
  assign multm_reduce_mc13 = multm_reduce_add3b0_maj3b_or3b_wx13 | multm_reduce_add3b0_maj3b_xy13;
  assign multm_reduce_mc14 = multm_reduce_add3b0_maj3b_or3b_wx14 | multm_reduce_add3b0_maj3b_xy14;
  assign multm_reduce_mc15 = multm_reduce_add3b0_maj3b_or3b_wx15 | multm_reduce_add3b0_maj3b_xy15;
  assign multm_reduce_mc16 = multm_reduce_add3b0_maj3b_or3b_wx16 | multm_reduce_add3b0_maj3b_xy16;
  assign multm_reduce_mc17 = multm_reduce_add3b0_maj3b_or3b_wx17 | multm_reduce_add3b0_maj3b_xy17;
  assign multm_reduce_mc18 = multm_reduce_add3b0_maj3b_or3b_wx18 | multm_reduce_add3b0_maj3b_xy18;
  assign multm_reduce_mc19 = multm_reduce_add3b0_maj3b_or3b_wx19 | multm_reduce_add3b0_maj3b_xy19;
  assign multm_reduce_mc20 = multm_reduce_add3b0_maj3b_or3b_wx20 | multm_reduce_add3b0_maj3b_xy20;
  assign multm_reduce_mc21 = multm_reduce_add3b0_maj3b_or3b_wx21 | multm_reduce_add3b0_maj3b_xy21;
  assign multm_reduce_mc22 = multm_reduce_add3b0_maj3b_or3b_wx22 | multm_reduce_add3b0_maj3b_xy22;
  assign multm_reduce_mc23 = multm_reduce_add3b0_maj3b_or3b_wx23 | multm_reduce_add3b0_maj3b_xy23;
  assign multm_reduce_mc24 = multm_reduce_add3b0_maj3b_or3b_wx24 | multm_reduce_add3b0_maj3b_xy24;
  assign multm_reduce_mc25 = multm_reduce_add3b0_maj3b_or3b_wx25 | multm_reduce_add3b0_maj3b_xy25;
  assign multm_reduce_mc26 = multm_reduce_add3b0_maj3b_or3b_wx26 | multm_reduce_add3b0_maj3b_xy26;
  assign multm_reduce_mc27 = multm_reduce_add3b0_maj3b_or3b_wx27 | multm_reduce_add3b0_maj3b_xy27;
  assign multm_reduce_mc28 = multm_reduce_add3b0_maj3b_or3b_wx28 | multm_reduce_add3b0_maj3b_xy28;
  assign multm_reduce_mc29 = multm_reduce_add3b0_maj3b_or3b_wx29 | multm_reduce_add3b0_maj3b_xy29;
  assign multm_reduce_mc30 = multm_reduce_add3b0_maj3b_or3b_wx30 | multm_reduce_add3b0_maj3b_xy30;
  assign multm_reduce_mc31 = multm_reduce_add3b0_maj3b_or3b_wx31 | multm_reduce_add3b0_maj3b_xy31;
  assign multm_reduce_mc32 = multm_reduce_add3b0_maj3b_or3b_wx32 | multm_reduce_add3b0_maj3b_xy32;
  assign multm_reduce_mc33 = multm_reduce_add3b0_maj3b_or3b_wx33 | multm_reduce_add3b0_maj3b_xy33;
  assign multm_reduce_mc34 = multm_reduce_add3b0_maj3b_or3b_wx34 | multm_reduce_add3b0_maj3b_xy34;
  assign multm_reduce_mc35 = multm_reduce_add3b0_maj3b_or3b_wx35 | multm_reduce_add3b0_maj3b_xy35;
  assign multm_reduce_mc36 = multm_reduce_add3b0_maj3b_or3b_wx36 | multm_reduce_add3b0_maj3b_xy36;
  assign multm_reduce_mc37 = multm_reduce_add3b0_maj3b_or3b_wx37 | multm_reduce_add3b0_maj3b_xy37;
  assign multm_reduce_mc38 = multm_reduce_add3b0_maj3b_or3b_wx38 | multm_reduce_add3b0_maj3b_xy38;
  assign multm_reduce_mc39 = multm_reduce_add3b0_maj3b_or3b_wx39 | multm_reduce_add3b0_maj3b_xy39;
  assign multm_reduce_mc40 = multm_reduce_add3b0_maj3b_or3b_wx40 | multm_reduce_add3b0_maj3b_xy40;
  assign multm_reduce_mc41 = multm_reduce_add3b0_maj3b_or3b_wx41 | multm_reduce_add3b0_maj3b_xy41;
  assign multm_reduce_mc42 = multm_reduce_add3b0_maj3b_or3b_wx42 | multm_reduce_add3b0_maj3b_xy42;
  assign multm_reduce_mc43 = multm_reduce_add3b0_maj3b_or3b_wx43 | multm_reduce_add3b0_maj3b_xy43;
  assign multm_reduce_mc44 = multm_reduce_add3b0_maj3b_or3b_wx44 | multm_reduce_add3b0_maj3b_xy44;
  assign multm_reduce_mc45 = multm_reduce_add3b0_maj3b_or3b_wx45 | multm_reduce_add3b0_maj3b_xy45;
  assign multm_reduce_mc46 = multm_reduce_add3b0_maj3b_or3b_wx46 | multm_reduce_add3b0_maj3b_xy46;
  assign multm_reduce_mc47 = multm_reduce_add3b0_maj3b_or3b_wx47 | multm_reduce_add3b0_maj3b_xy47;
  assign multm_reduce_mc48 = multm_reduce_add3b0_maj3b_or3b_wx48 | multm_reduce_add3b0_maj3b_xy48;
  assign multm_reduce_mc49 = multm_reduce_add3b0_maj3b_or3b_wx49 | multm_reduce_add3b0_maj3b_xy49;
  assign multm_reduce_mc50 = multm_reduce_add3b0_maj3b_or3b_wx50 | multm_reduce_add3b0_maj3b_xy50;
  assign multm_reduce_mc51 = multm_reduce_add3b0_maj3b_or3b_wx51 | multm_reduce_add3b0_maj3b_xy51;
  assign multm_reduce_mc52 = multm_reduce_add3b0_maj3b_or3b_wx52 | multm_reduce_add3b0_maj3b_xy52;
  assign multm_reduce_mc53 = multm_reduce_add3b0_maj3b_or3b_wx53 | multm_reduce_add3b0_maj3b_xy53;
  assign multm_reduce_mc54 = multm_reduce_add3b0_maj3b_or3b_wx54 | multm_reduce_add3b0_maj3b_xy54;
  assign multm_reduce_mc55 = multm_reduce_add3b0_maj3b_or3b_wx55 | multm_reduce_add3b0_maj3b_xy55;
  assign multm_reduce_mc56 = multm_reduce_add3b0_maj3b_or3b_wx56 | multm_reduce_add3b0_maj3b_xy56;
  assign multm_reduce_mc57 = multm_reduce_add3b0_maj3b_or3b_wx57 | multm_reduce_add3b0_maj3b_xy57;
  assign multm_reduce_mc58 = multm_reduce_add3b0_maj3b_or3b_wx58 | multm_reduce_add3b0_maj3b_xy58;
  assign multm_reduce_mc59 = multm_reduce_add3b0_maj3b_or3b_wx59 | multm_reduce_add3b0_maj3b_xy59;
  assign multm_reduce_mc60 = multm_reduce_add3b0_maj3b_or3b_wx60 | multm_reduce_add3b0_maj3b_xy60;
  assign multm_reduce_mc61 = multm_reduce_add3b0_maj3b_or3b_wx61 | multm_reduce_add3b0_maj3b_xy61;
  assign multm_reduce_mc62 = multm_reduce_add3b0_maj3b_or3b_wx62 | multm_reduce_add3b0_maj3b_xy62;
  assign multm_reduce_mc63 = multm_reduce_add3b0_maj3b_or3b_wx63 | multm_reduce_add3b0_maj3b_xy63;
  assign multm_reduce_mc64 = multm_reduce_add3b0_maj3b_or3b_wx64 | multm_reduce_add3b0_maj3b_xy64;
  assign multm_reduce_mc65 = multm_reduce_add3b0_maj3b_or3b_wx65 | multm_reduce_add3b0_maj3b_xy65;
  assign multm_reduce_mc66 = multm_reduce_add3b0_maj3b_or3b_wx66 | multm_reduce_add3b0_maj3b_xy66;
  assign multm_reduce_mc67 = multm_reduce_add3b0_maj3b_or3b_wx67 | multm_reduce_add3b0_maj3b_xy67;
  assign multm_reduce_mc68 = multm_reduce_add3b0_maj3b_or3b_wx68 | multm_reduce_add3b0_maj3b_xy68;
  assign multm_reduce_mc69 = multm_reduce_add3b0_maj3b_or3b_wx69 | multm_reduce_add3b0_maj3b_xy69;
  assign multm_reduce_mc70 = multm_reduce_add3b0_maj3b_or3b_wx70 | multm_reduce_add3b0_maj3b_xy70;
  assign multm_reduce_mc71 = multm_reduce_add3b0_maj3b_or3b_wx71 | multm_reduce_add3b0_maj3b_xy71;
  assign multm_reduce_mc72 = multm_reduce_add3b0_maj3b_or3b_wx72 | multm_reduce_add3b0_maj3b_xy72;
  assign multm_reduce_mc73 = multm_reduce_add3b0_maj3b_or3b_wx73 | multm_reduce_add3b0_maj3b_xy73;
  assign multm_reduce_mc74 = multm_reduce_add3b0_maj3b_or3b_wx74 | multm_reduce_add3b0_maj3b_xy74;
  assign multm_reduce_mc75 = multm_reduce_add3b0_maj3b_or3b_wx75 | multm_reduce_add3b0_maj3b_xy75;
  assign multm_reduce_mc76 = multm_reduce_add3b0_maj3b_or3b_wx76 | multm_reduce_add3b0_maj3b_xy76;
  assign multm_reduce_mc77 = multm_reduce_add3b0_maj3b_or3b_wx77 | multm_reduce_add3b0_maj3b_xy77;
  assign multm_reduce_mc78 = multm_reduce_add3b0_maj3b_or3b_wx78 | multm_reduce_add3b0_maj3b_xy78;
  assign multm_reduce_mc79 = multm_reduce_add3b0_maj3b_or3b_wx79 | multm_reduce_add3b0_maj3b_xy79;
  assign multm_reduce_mc80 = multm_reduce_add3b0_maj3b_or3b_wx80 | multm_reduce_add3b0_maj3b_xy80;
  assign multm_reduce_mc81 = multm_reduce_add3b0_maj3b_or3b_wx81 | multm_reduce_add3b0_maj3b_xy81;
  assign multm_reduce_mc82 = multm_reduce_add3b0_maj3b_or3b_wx82 | multm_reduce_add3b0_maj3b_xy82;
  assign multm_reduce_mc83 = multm_reduce_add3b0_maj3b_or3b_wx83 | multm_reduce_add3b0_maj3b_xy83;
  assign multm_reduce_mc84 = multm_reduce_add3b0_maj3b_or3b_wx84 | multm_reduce_add3b0_maj3b_xy84;
  assign multm_reduce_mc85 = multm_reduce_add3b0_maj3b_or3b_wx85 | multm_reduce_add3b0_maj3b_xy85;
  assign multm_reduce_mc86 = multm_reduce_add3b0_maj3b_or3b_wx86 | multm_reduce_add3b0_maj3b_xy86;
  assign multm_reduce_mc87 = multm_reduce_add3b0_maj3b_or3b_wx87 | multm_reduce_add3b0_maj3b_xy87;
  assign multm_reduce_mc88 = multm_reduce_add3b0_maj3b_or3b_wx88 | multm_reduce_add3b0_maj3b_xy88;
  assign multm_reduce_mc89 = multm_reduce_add3b0_maj3b_or3b_wx89 | multm_reduce_add3b0_maj3b_xy89;
  assign multm_reduce_mc90 = multm_reduce_add3b0_maj3b_or3b_wx90 | multm_reduce_add3b0_maj3b_xy90;
  assign multm_reduce_mc91 = multm_reduce_add3b0_maj3b_or3b_wx91 | multm_reduce_add3b0_maj3b_xy91;
  assign multm_reduce_mc92 = multm_reduce_add3b0_maj3b_or3b_wx92 | multm_reduce_add3b0_maj3b_xy92;
  assign multm_reduce_mc93 = multm_reduce_add3b0_maj3b_or3b_wx93 | multm_reduce_add3b0_maj3b_xy93;
  assign multm_reduce_mc94 = multm_reduce_add3b0_maj3b_or3b_wx94 | multm_reduce_add3b0_maj3b_xy94;
  assign multm_reduce_mc95 = multm_reduce_add3b0_maj3b_or3b_wx95 | multm_reduce_add3b0_maj3b_xy95;
  assign multm_reduce_mc96 = multm_reduce_add3b0_maj3b_or3b_wx96 | multm_reduce_add3b0_maj3b_xy96;
  assign multm_reduce_mc97 = multm_reduce_add3b0_maj3b_or3b_wx97 | multm_reduce_add3b0_maj3b_xy97;
  assign multm_reduce_mc98 = multm_reduce_add3b0_maj3b_or3b_wx98 | multm_reduce_add3b0_maj3b_xy98;
  assign multm_reduce_mc99 = multm_reduce_add3b0_maj3b_or3b_wx99 | multm_reduce_add3b0_maj3b_xy99;
  assign multm_reduce_mc100 = multm_reduce_add3b0_maj3b_or3b_wx100 | multm_reduce_add3b0_maj3b_xy100;
  assign multm_reduce_mc101 = multm_reduce_add3b0_maj3b_or3b_wx101 | multm_reduce_add3b0_maj3b_xy101;
  assign multm_reduce_mc102 = multm_reduce_add3b0_maj3b_or3b_wx102 | multm_reduce_add3b0_maj3b_xy102;
  assign multm_reduce_mc103 = multm_reduce_add3b0_maj3b_or3b_wx103 | multm_reduce_add3b0_maj3b_xy103;
  assign multm_reduce_mc104 = multm_reduce_add3b0_maj3b_or3b_wx104 | multm_reduce_add3b0_maj3b_xy104;
  assign multm_reduce_mc105 = multm_reduce_add3b0_maj3b_or3b_wx105 | multm_reduce_add3b0_maj3b_xy105;
  assign multm_reduce_mc106 = multm_reduce_add3b0_maj3b_or3b_wx106 | multm_reduce_add3b0_maj3b_xy106;
  assign multm_reduce_mc107 = multm_reduce_add3b0_maj3b_or3b_wx107 | multm_reduce_add3b0_maj3b_xy107;
  assign multm_reduce_mc108 = multm_reduce_add3b0_maj3b_or3b_wx108 | multm_reduce_add3b0_maj3b_xy108;
  assign multm_reduce_mc109 = multm_reduce_add3b0_maj3b_or3b_wx109 | multm_reduce_add3b0_maj3b_xy109;
  assign multm_reduce_mc110 = multm_reduce_add3b0_maj3b_or3b_wx110 | multm_reduce_add3b0_maj3b_xy110;
  assign multm_reduce_mc111 = multm_reduce_add3b0_maj3b_or3b_wx111 | multm_reduce_add3b0_maj3b_xy111;
  assign multm_reduce_mc112 = multm_reduce_add3b0_maj3b_or3b_wx112 | multm_reduce_add3b0_maj3b_xy112;
  assign multm_reduce_mc113 = multm_reduce_add3b0_maj3b_or3b_wx113 | multm_reduce_add3b0_maj3b_xy113;
  assign multm_reduce_mc114 = multm_reduce_add3b0_maj3b_or3b_wx114 | multm_reduce_add3b0_maj3b_xy114;
  assign multm_reduce_mc115 = multm_reduce_add3b0_maj3b_or3b_wx115 | multm_reduce_add3b0_maj3b_xy115;
  assign multm_reduce_mc116 = multm_reduce_add3b0_maj3b_or3b_wx116 | multm_reduce_add3b0_maj3b_xy116;
  assign multm_reduce_mc117 = multm_reduce_add3b0_maj3b_or3b_wx117 | multm_reduce_add3b0_maj3b_xy117;
  assign multm_reduce_mc118 = multm_reduce_add3b0_maj3b_or3b_wx118 | multm_reduce_add3b0_maj3b_xy118;
  assign multm_reduce_mc119 = multm_reduce_add3b0_maj3b_or3b_wx119 | multm_reduce_add3b0_maj3b_xy119;
  assign multm_reduce_mc120 = multm_reduce_add3b0_maj3b_or3b_wx120 | multm_reduce_add3b0_maj3b_xy120;
  assign multm_reduce_mc121 = multm_reduce_add3b0_maj3b_or3b_wx121 | multm_reduce_add3b0_maj3b_xy121;
  assign multm_reduce_mc122 = multm_reduce_add3b0_maj3b_or3b_wx122 | multm_reduce_add3b0_maj3b_xy122;
  assign multm_reduce_mc123 = multm_reduce_add3b0_maj3b_or3b_wx123 | multm_reduce_add3b0_maj3b_xy123;
  assign multm_reduce_mc124 = multm_reduce_add3b0_maj3b_or3b_wx124 | multm_reduce_add3b0_maj3b_xy124;
  assign multm_reduce_mc125 = multm_reduce_add3b0_maj3b_or3b_wx125 | multm_reduce_add3b0_maj3b_xy125;
  assign multm_reduce_mc126 = multm_reduce_add3b0_maj3b_or3b_wx126 | multm_reduce_add3b0_maj3b_xy126;
  assign multm_reduce_mc127 = multm_reduce_add3b0_maj3b_or3b_wx127 | multm_reduce_add3b0_maj3b_xy127;
  assign multm_reduce_mc128 = multm_reduce_add3b0_maj3b_or3b_wx128 | multm_reduce_add3b0_maj3b_xy128;
  assign multm_reduce_mc129 = multm_reduce_add3b0_maj3b_or3b_wx129 | multm_reduce_add3b0_maj3b_xy129;
  assign multm_reduce_mc130 = multm_reduce_add3b0_maj3b_or3b_wx130 | multm_reduce_add3b0_maj3b_xy130;
  assign multm_reduce_mc131 = multm_reduce_add3b0_maj3b_or3b_wx131 | multm_reduce_add3b0_maj3b_xy131;
  assign multm_reduce_mc132 = multm_reduce_add3b0_maj3b_or3b_wx132 | multm_reduce_add3b0_maj3b_xy132;
  assign multm_reduce_mc133 = multm_reduce_add3b0_maj3b_or3b_wx133 | multm_reduce_add3b0_maj3b_xy133;
  assign multm_reduce_mc134 = multm_reduce_add3b0_maj3b_or3b_wx134 | multm_reduce_add3b0_maj3b_xy134;
  assign multm_reduce_mc135 = multm_reduce_add3b0_maj3b_or3b_wx135 | multm_reduce_add3b0_maj3b_xy135;
  assign multm_reduce_mc136 = multm_reduce_add3b0_maj3b_or3b_wx136 | multm_reduce_add3b0_maj3b_xy136;
  assign multm_reduce_mc137 = multm_reduce_add3b0_maj3b_or3b_wx137 | multm_reduce_add3b0_maj3b_xy137;
  assign multm_reduce_mc138 = multm_reduce_add3b0_maj3b_or3b_wx138 | multm_reduce_add3b0_maj3b_xy138;
  assign multm_reduce_mc139 = multm_reduce_add3b0_maj3b_or3b_wx139 | multm_reduce_add3b0_maj3b_xy139;
  assign multm_reduce_mc140 = multm_reduce_add3b0_maj3b_or3b_wx140 | multm_reduce_add3b0_maj3b_xy140;
  assign multm_reduce_mc141 = multm_reduce_add3b0_maj3b_or3b_wx141 | multm_reduce_add3b0_maj3b_xy141;
  assign multm_reduce_mc142 = multm_reduce_add3b0_maj3b_or3b_wx142 | multm_reduce_add3b0_maj3b_xy142;
  assign multm_reduce_mc143 = multm_reduce_add3b0_maj3b_or3b_wx143 | multm_reduce_add3b0_maj3b_xy143;
  assign multm_reduce_mc144 = multm_reduce_add3b0_maj3b_or3b_wx144 | multm_reduce_add3b0_maj3b_xy144;
  assign multm_reduce_mc145 = multm_reduce_add3b0_maj3b_or3b_wx145 | multm_reduce_add3b0_maj3b_xy145;
  assign multm_reduce_mc146 = multm_reduce_add3b0_maj3b_or3b_wx146 | multm_reduce_add3b0_maj3b_xy146;
  assign multm_reduce_mc147 = multm_reduce_add3b0_maj3b_or3b_wx147 | multm_reduce_add3b0_maj3b_xy147;
  assign multm_reduce_mc148 = multm_reduce_add3b0_maj3b_or3b_wx148 | multm_reduce_add3b0_maj3b_xy148;
  assign multm_reduce_mc149 = multm_reduce_add3b0_maj3b_or3b_wx149 | multm_reduce_add3b0_maj3b_xy149;
  assign multm_reduce_mc150 = multm_reduce_add3b0_maj3b_or3b_wx150 | multm_reduce_add3b0_maj3b_xy150;
  assign multm_reduce_mc151 = multm_reduce_add3b0_maj3b_or3b_wx151 | multm_reduce_add3b0_maj3b_xy151;
  assign multm_reduce_mc152 = multm_reduce_add3b0_maj3b_or3b_wx152 | multm_reduce_add3b0_maj3b_xy152;
  assign multm_reduce_mc153 = multm_reduce_add3b0_maj3b_or3b_wx153 | multm_reduce_add3b0_maj3b_xy153;
  assign multm_reduce_mc154 = multm_reduce_add3b0_maj3b_or3b_wx154 | multm_reduce_add3b0_maj3b_xy154;
  assign multm_reduce_mc155 = multm_reduce_add3b0_maj3b_or3b_wx155 | multm_reduce_add3b0_maj3b_xy155;
  assign multm_reduce_mc156 = multm_reduce_add3b0_maj3b_or3b_wx156 | multm_reduce_add3b0_maj3b_xy156;
  assign multm_reduce_mc157 = multm_reduce_add3b0_maj3b_or3b_wx157 | multm_reduce_add3b0_maj3b_xy157;
  assign multm_reduce_mc158 = multm_reduce_add3b0_maj3b_or3b_wx158 | multm_reduce_add3b0_maj3b_xy158;
  assign multm_reduce_mc159 = multm_reduce_add3b0_maj3b_or3b_wx159 | multm_reduce_add3b0_maj3b_xy159;
  assign multm_reduce_mc160 = multm_reduce_add3b0_maj3b_or3b_wx160 | multm_reduce_add3b0_maj3b_xy160;
  assign multm_reduce_mc161 = multm_reduce_add3b0_maj3b_or3b_wx161 | multm_reduce_add3b0_maj3b_xy161;
  assign multm_reduce_mc162 = multm_reduce_add3b0_maj3b_or3b_wx162 | multm_reduce_add3b0_maj3b_xy162;
  assign multm_reduce_mc163 = multm_reduce_add3b0_maj3b_or3b_wx163 | multm_reduce_add3b0_maj3b_xy163;
  assign multm_reduce_mc164 = multm_reduce_add3b0_maj3b_or3b_wx164 | multm_reduce_add3b0_maj3b_xy164;
  assign multm_reduce_mc165 = multm_reduce_add3b0_maj3b_or3b_wx165 | multm_reduce_add3b0_maj3b_xy165;
  assign multm_reduce_mc166 = multm_reduce_add3b0_maj3b_or3b_wx166 | multm_reduce_add3b0_maj3b_xy166;
  assign multm_reduce_mc167 = multm_reduce_add3b0_maj3b_or3b_wx167 | multm_reduce_add3b0_maj3b_xy167;
  assign multm_reduce_mc168 = multm_reduce_add3b0_maj3b_or3b_wx168 | multm_reduce_add3b0_maj3b_xy168;
  assign multm_reduce_mc169 = multm_reduce_add3b0_maj3b_or3b_wx169 | multm_reduce_add3b0_maj3b_xy169;
  assign multm_reduce_mc170 = multm_reduce_add3b0_maj3b_or3b_wx170 | multm_reduce_add3b0_maj3b_xy170;
  assign multm_reduce_mc171 = multm_reduce_add3b0_maj3b_or3b_wx171 | multm_reduce_add3b0_maj3b_xy171;
  assign multm_reduce_mc172 = multm_reduce_add3b0_maj3b_or3b_wx172 | multm_reduce_add3b0_maj3b_xy172;
  assign multm_reduce_mc173 = multm_reduce_add3b0_maj3b_or3b_wx173 | multm_reduce_add3b0_maj3b_xy173;
  assign multm_reduce_mc174 = multm_reduce_add3b0_maj3b_or3b_wx174 | multm_reduce_add3b0_maj3b_xy174;
  assign multm_reduce_mc175 = multm_reduce_add3b0_maj3b_or3b_wx175 | multm_reduce_add3b0_maj3b_xy175;
  assign multm_reduce_mc176 = multm_reduce_add3b0_maj3b_or3b_wx176 | multm_reduce_add3b0_maj3b_xy176;
  assign multm_reduce_mc177 = multm_reduce_add3b0_maj3b_or3b_wx177 | multm_reduce_add3b0_maj3b_xy177;
  assign multm_reduce_mc178 = multm_reduce_add3b0_maj3b_or3b_wx178 | multm_reduce_add3b0_maj3b_xy178;
  assign multm_reduce_mc179 = multm_reduce_add3b0_maj3b_or3b_wx179 | multm_reduce_add3b0_maj3b_xy179;
  assign multm_reduce_mc180 = multm_reduce_add3b0_maj3b_or3b_wx180 | multm_reduce_add3b0_maj3b_xy180;
  assign multm_reduce_mc181 = multm_reduce_add3b0_maj3b_or3b_wx181 | multm_reduce_add3b0_maj3b_xy181;
  assign multm_reduce_mc182 = multm_reduce_add3b0_maj3b_or3b_wx182 | multm_reduce_add3b0_maj3b_xy182;
  assign multm_reduce_mc183 = multm_reduce_sa183 & multm_reduce_sd183;
  assign multm_reduce_ms11 = multm_reduce_add3b0_xor3b_wx11 ^ multm_reduce_sd11;
  assign multm_reduce_ms12 = multm_reduce_add3b0_xor3b_wx12 ^ multm_reduce_sd12;
  assign multm_reduce_ms13 = multm_reduce_add3b0_xor3b_wx13 ^ multm_reduce_sd13;
  assign multm_reduce_ms14 = multm_reduce_add3b0_xor3b_wx14 ^ multm_reduce_sd14;
  assign multm_reduce_ms15 = multm_reduce_add3b0_xor3b_wx15 ^ multm_reduce_sd15;
  assign multm_reduce_ms16 = multm_reduce_add3b0_xor3b_wx16 ^ multm_reduce_sd16;
  assign multm_reduce_ms17 = multm_reduce_add3b0_xor3b_wx17 ^ multm_reduce_sd17;
  assign multm_reduce_ms18 = multm_reduce_add3b0_xor3b_wx18 ^ multm_reduce_sd18;
  assign multm_reduce_ms19 = multm_reduce_add3b0_xor3b_wx19 ^ multm_reduce_sd19;
  assign multm_reduce_ms20 = multm_reduce_add3b0_xor3b_wx20 ^ multm_reduce_sd20;
  assign multm_reduce_ms21 = multm_reduce_add3b0_xor3b_wx21 ^ multm_reduce_sd21;
  assign multm_reduce_ms22 = multm_reduce_add3b0_xor3b_wx22 ^ multm_reduce_sd22;
  assign multm_reduce_ms23 = multm_reduce_add3b0_xor3b_wx23 ^ multm_reduce_sd23;
  assign multm_reduce_ms24 = multm_reduce_add3b0_xor3b_wx24 ^ multm_reduce_sd24;
  assign multm_reduce_ms25 = multm_reduce_add3b0_xor3b_wx25 ^ multm_reduce_sd25;
  assign multm_reduce_ms26 = multm_reduce_add3b0_xor3b_wx26 ^ multm_reduce_sd26;
  assign multm_reduce_ms27 = multm_reduce_add3b0_xor3b_wx27 ^ multm_reduce_sd27;
  assign multm_reduce_ms28 = multm_reduce_add3b0_xor3b_wx28 ^ multm_reduce_sd28;
  assign multm_reduce_ms29 = multm_reduce_add3b0_xor3b_wx29 ^ multm_reduce_sd29;
  assign multm_reduce_ms30 = multm_reduce_add3b0_xor3b_wx30 ^ multm_reduce_sd30;
  assign multm_reduce_ms31 = multm_reduce_add3b0_xor3b_wx31 ^ multm_reduce_sd31;
  assign multm_reduce_ms32 = multm_reduce_add3b0_xor3b_wx32 ^ multm_reduce_sd32;
  assign multm_reduce_ms33 = multm_reduce_add3b0_xor3b_wx33 ^ multm_reduce_sd33;
  assign multm_reduce_ms34 = multm_reduce_add3b0_xor3b_wx34 ^ multm_reduce_sd34;
  assign multm_reduce_ms35 = multm_reduce_add3b0_xor3b_wx35 ^ multm_reduce_sd35;
  assign multm_reduce_ms36 = multm_reduce_add3b0_xor3b_wx36 ^ multm_reduce_sd36;
  assign multm_reduce_ms37 = multm_reduce_add3b0_xor3b_wx37 ^ multm_reduce_sd37;
  assign multm_reduce_ms38 = multm_reduce_add3b0_xor3b_wx38 ^ multm_reduce_sd38;
  assign multm_reduce_ms39 = multm_reduce_add3b0_xor3b_wx39 ^ multm_reduce_sd39;
  assign multm_reduce_ms40 = multm_reduce_add3b0_xor3b_wx40 ^ multm_reduce_sd40;
  assign multm_reduce_ms41 = multm_reduce_add3b0_xor3b_wx41 ^ multm_reduce_sd41;
  assign multm_reduce_ms42 = multm_reduce_add3b0_xor3b_wx42 ^ multm_reduce_sd42;
  assign multm_reduce_ms43 = multm_reduce_add3b0_xor3b_wx43 ^ multm_reduce_sd43;
  assign multm_reduce_ms44 = multm_reduce_add3b0_xor3b_wx44 ^ multm_reduce_sd44;
  assign multm_reduce_ms45 = multm_reduce_add3b0_xor3b_wx45 ^ multm_reduce_sd45;
  assign multm_reduce_ms46 = multm_reduce_add3b0_xor3b_wx46 ^ multm_reduce_sd46;
  assign multm_reduce_ms47 = multm_reduce_add3b0_xor3b_wx47 ^ multm_reduce_sd47;
  assign multm_reduce_ms48 = multm_reduce_add3b0_xor3b_wx48 ^ multm_reduce_sd48;
  assign multm_reduce_ms49 = multm_reduce_add3b0_xor3b_wx49 ^ multm_reduce_sd49;
  assign multm_reduce_ms50 = multm_reduce_add3b0_xor3b_wx50 ^ multm_reduce_sd50;
  assign multm_reduce_ms51 = multm_reduce_add3b0_xor3b_wx51 ^ multm_reduce_sd51;
  assign multm_reduce_ms52 = multm_reduce_add3b0_xor3b_wx52 ^ multm_reduce_sd52;
  assign multm_reduce_ms53 = multm_reduce_add3b0_xor3b_wx53 ^ multm_reduce_sd53;
  assign multm_reduce_ms54 = multm_reduce_add3b0_xor3b_wx54 ^ multm_reduce_sd54;
  assign multm_reduce_ms55 = multm_reduce_add3b0_xor3b_wx55 ^ multm_reduce_sd55;
  assign multm_reduce_ms56 = multm_reduce_add3b0_xor3b_wx56 ^ multm_reduce_sd56;
  assign multm_reduce_ms57 = multm_reduce_add3b0_xor3b_wx57 ^ multm_reduce_sd57;
  assign multm_reduce_ms58 = multm_reduce_add3b0_xor3b_wx58 ^ multm_reduce_sd58;
  assign multm_reduce_ms59 = multm_reduce_add3b0_xor3b_wx59 ^ multm_reduce_sd59;
  assign multm_reduce_ms60 = multm_reduce_add3b0_xor3b_wx60 ^ multm_reduce_sd60;
  assign multm_reduce_ms61 = multm_reduce_add3b0_xor3b_wx61 ^ multm_reduce_sd61;
  assign multm_reduce_ms62 = multm_reduce_add3b0_xor3b_wx62 ^ multm_reduce_sd62;
  assign multm_reduce_ms63 = multm_reduce_add3b0_xor3b_wx63 ^ multm_reduce_sd63;
  assign multm_reduce_ms64 = multm_reduce_add3b0_xor3b_wx64 ^ multm_reduce_sd64;
  assign multm_reduce_ms65 = multm_reduce_add3b0_xor3b_wx65 ^ multm_reduce_sd65;
  assign multm_reduce_ms66 = multm_reduce_add3b0_xor3b_wx66 ^ multm_reduce_sd66;
  assign multm_reduce_ms67 = multm_reduce_add3b0_xor3b_wx67 ^ multm_reduce_sd67;
  assign multm_reduce_ms68 = multm_reduce_add3b0_xor3b_wx68 ^ multm_reduce_sd68;
  assign multm_reduce_ms69 = multm_reduce_add3b0_xor3b_wx69 ^ multm_reduce_sd69;
  assign multm_reduce_ms70 = multm_reduce_add3b0_xor3b_wx70 ^ multm_reduce_sd70;
  assign multm_reduce_ms71 = multm_reduce_add3b0_xor3b_wx71 ^ multm_reduce_sd71;
  assign multm_reduce_ms72 = multm_reduce_add3b0_xor3b_wx72 ^ multm_reduce_sd72;
  assign multm_reduce_ms73 = multm_reduce_add3b0_xor3b_wx73 ^ multm_reduce_sd73;
  assign multm_reduce_ms74 = multm_reduce_add3b0_xor3b_wx74 ^ multm_reduce_sd74;
  assign multm_reduce_ms75 = multm_reduce_add3b0_xor3b_wx75 ^ multm_reduce_sd75;
  assign multm_reduce_ms76 = multm_reduce_add3b0_xor3b_wx76 ^ multm_reduce_sd76;
  assign multm_reduce_ms77 = multm_reduce_add3b0_xor3b_wx77 ^ multm_reduce_sd77;
  assign multm_reduce_ms78 = multm_reduce_add3b0_xor3b_wx78 ^ multm_reduce_sd78;
  assign multm_reduce_ms79 = multm_reduce_add3b0_xor3b_wx79 ^ multm_reduce_sd79;
  assign multm_reduce_ms80 = multm_reduce_add3b0_xor3b_wx80 ^ multm_reduce_sd80;
  assign multm_reduce_ms81 = multm_reduce_add3b0_xor3b_wx81 ^ multm_reduce_sd81;
  assign multm_reduce_ms82 = multm_reduce_add3b0_xor3b_wx82 ^ multm_reduce_sd82;
  assign multm_reduce_ms83 = multm_reduce_add3b0_xor3b_wx83 ^ multm_reduce_sd83;
  assign multm_reduce_ms84 = multm_reduce_add3b0_xor3b_wx84 ^ multm_reduce_sd84;
  assign multm_reduce_ms85 = multm_reduce_add3b0_xor3b_wx85 ^ multm_reduce_sd85;
  assign multm_reduce_ms86 = multm_reduce_add3b0_xor3b_wx86 ^ multm_reduce_sd86;
  assign multm_reduce_ms87 = multm_reduce_add3b0_xor3b_wx87 ^ multm_reduce_sd87;
  assign multm_reduce_ms88 = multm_reduce_add3b0_xor3b_wx88 ^ multm_reduce_sd88;
  assign multm_reduce_ms89 = multm_reduce_add3b0_xor3b_wx89 ^ multm_reduce_sd89;
  assign multm_reduce_ms90 = multm_reduce_add3b0_xor3b_wx90 ^ multm_reduce_sd90;
  assign multm_reduce_ms91 = multm_reduce_add3b0_xor3b_wx91 ^ multm_reduce_sd91;
  assign multm_reduce_ms92 = multm_reduce_add3b0_xor3b_wx92 ^ multm_reduce_sd92;
  assign multm_reduce_ms93 = multm_reduce_add3b0_xor3b_wx93 ^ multm_reduce_sd93;
  assign multm_reduce_ms94 = multm_reduce_add3b0_xor3b_wx94 ^ multm_reduce_sd94;
  assign multm_reduce_ms95 = multm_reduce_add3b0_xor3b_wx95 ^ multm_reduce_sd95;
  assign multm_reduce_ms96 = multm_reduce_add3b0_xor3b_wx96 ^ multm_reduce_sd96;
  assign multm_reduce_ms97 = multm_reduce_add3b0_xor3b_wx97 ^ multm_reduce_sd97;
  assign multm_reduce_ms98 = multm_reduce_add3b0_xor3b_wx98 ^ multm_reduce_sd98;
  assign multm_reduce_ms99 = multm_reduce_add3b0_xor3b_wx99 ^ multm_reduce_sd99;
  assign multm_reduce_ms100 = multm_reduce_add3b0_xor3b_wx100 ^ multm_reduce_sd100;
  assign multm_reduce_ms101 = multm_reduce_add3b0_xor3b_wx101 ^ multm_reduce_sd101;
  assign multm_reduce_ms102 = multm_reduce_add3b0_xor3b_wx102 ^ multm_reduce_sd102;
  assign multm_reduce_ms103 = multm_reduce_add3b0_xor3b_wx103 ^ multm_reduce_sd103;
  assign multm_reduce_ms104 = multm_reduce_add3b0_xor3b_wx104 ^ multm_reduce_sd104;
  assign multm_reduce_ms105 = multm_reduce_add3b0_xor3b_wx105 ^ multm_reduce_sd105;
  assign multm_reduce_ms106 = multm_reduce_add3b0_xor3b_wx106 ^ multm_reduce_sd106;
  assign multm_reduce_ms107 = multm_reduce_add3b0_xor3b_wx107 ^ multm_reduce_sd107;
  assign multm_reduce_ms108 = multm_reduce_add3b0_xor3b_wx108 ^ multm_reduce_sd108;
  assign multm_reduce_ms109 = multm_reduce_add3b0_xor3b_wx109 ^ multm_reduce_sd109;
  assign multm_reduce_ms110 = multm_reduce_add3b0_xor3b_wx110 ^ multm_reduce_sd110;
  assign multm_reduce_ms111 = multm_reduce_add3b0_xor3b_wx111 ^ multm_reduce_sd111;
  assign multm_reduce_ms112 = multm_reduce_add3b0_xor3b_wx112 ^ multm_reduce_sd112;
  assign multm_reduce_ms113 = multm_reduce_add3b0_xor3b_wx113 ^ multm_reduce_sd113;
  assign multm_reduce_ms114 = multm_reduce_add3b0_xor3b_wx114 ^ multm_reduce_sd114;
  assign multm_reduce_ms115 = multm_reduce_add3b0_xor3b_wx115 ^ multm_reduce_sd115;
  assign multm_reduce_ms116 = multm_reduce_add3b0_xor3b_wx116 ^ multm_reduce_sd116;
  assign multm_reduce_ms117 = multm_reduce_add3b0_xor3b_wx117 ^ multm_reduce_sd117;
  assign multm_reduce_ms118 = multm_reduce_add3b0_xor3b_wx118 ^ multm_reduce_sd118;
  assign multm_reduce_ms119 = multm_reduce_add3b0_xor3b_wx119 ^ multm_reduce_sd119;
  assign multm_reduce_ms120 = multm_reduce_add3b0_xor3b_wx120 ^ multm_reduce_sd120;
  assign multm_reduce_ms121 = multm_reduce_add3b0_xor3b_wx121 ^ multm_reduce_sd121;
  assign multm_reduce_ms122 = multm_reduce_add3b0_xor3b_wx122 ^ multm_reduce_sd122;
  assign multm_reduce_ms123 = multm_reduce_add3b0_xor3b_wx123 ^ multm_reduce_sd123;
  assign multm_reduce_ms124 = multm_reduce_add3b0_xor3b_wx124 ^ multm_reduce_sd124;
  assign multm_reduce_ms125 = multm_reduce_add3b0_xor3b_wx125 ^ multm_reduce_sd125;
  assign multm_reduce_ms126 = multm_reduce_add3b0_xor3b_wx126 ^ multm_reduce_sd126;
  assign multm_reduce_ms127 = multm_reduce_add3b0_xor3b_wx127 ^ multm_reduce_sd127;
  assign multm_reduce_ms128 = multm_reduce_add3b0_xor3b_wx128 ^ multm_reduce_sd128;
  assign multm_reduce_ms129 = multm_reduce_add3b0_xor3b_wx129 ^ multm_reduce_sd129;
  assign multm_reduce_ms130 = multm_reduce_add3b0_xor3b_wx130 ^ multm_reduce_sd130;
  assign multm_reduce_ms131 = multm_reduce_add3b0_xor3b_wx131 ^ multm_reduce_sd131;
  assign multm_reduce_ms132 = multm_reduce_add3b0_xor3b_wx132 ^ multm_reduce_sd132;
  assign multm_reduce_ms133 = multm_reduce_add3b0_xor3b_wx133 ^ multm_reduce_sd133;
  assign multm_reduce_ms134 = multm_reduce_add3b0_xor3b_wx134 ^ multm_reduce_sd134;
  assign multm_reduce_ms135 = multm_reduce_add3b0_xor3b_wx135 ^ multm_reduce_sd135;
  assign multm_reduce_ms136 = multm_reduce_add3b0_xor3b_wx136 ^ multm_reduce_sd136;
  assign multm_reduce_ms137 = multm_reduce_add3b0_xor3b_wx137 ^ multm_reduce_sd137;
  assign multm_reduce_ms138 = multm_reduce_add3b0_xor3b_wx138 ^ multm_reduce_sd138;
  assign multm_reduce_ms139 = multm_reduce_add3b0_xor3b_wx139 ^ multm_reduce_sd139;
  assign multm_reduce_ms140 = multm_reduce_add3b0_xor3b_wx140 ^ multm_reduce_sd140;
  assign multm_reduce_ms141 = multm_reduce_add3b0_xor3b_wx141 ^ multm_reduce_sd141;
  assign multm_reduce_ms142 = multm_reduce_add3b0_xor3b_wx142 ^ multm_reduce_sd142;
  assign multm_reduce_ms143 = multm_reduce_add3b0_xor3b_wx143 ^ multm_reduce_sd143;
  assign multm_reduce_ms144 = multm_reduce_add3b0_xor3b_wx144 ^ multm_reduce_sd144;
  assign multm_reduce_ms145 = multm_reduce_add3b0_xor3b_wx145 ^ multm_reduce_sd145;
  assign multm_reduce_ms146 = multm_reduce_add3b0_xor3b_wx146 ^ multm_reduce_sd146;
  assign multm_reduce_ms147 = multm_reduce_add3b0_xor3b_wx147 ^ multm_reduce_sd147;
  assign multm_reduce_ms148 = multm_reduce_add3b0_xor3b_wx148 ^ multm_reduce_sd148;
  assign multm_reduce_ms149 = multm_reduce_add3b0_xor3b_wx149 ^ multm_reduce_sd149;
  assign multm_reduce_ms150 = multm_reduce_add3b0_xor3b_wx150 ^ multm_reduce_sd150;
  assign multm_reduce_ms151 = multm_reduce_add3b0_xor3b_wx151 ^ multm_reduce_sd151;
  assign multm_reduce_ms152 = multm_reduce_add3b0_xor3b_wx152 ^ multm_reduce_sd152;
  assign multm_reduce_ms153 = multm_reduce_add3b0_xor3b_wx153 ^ multm_reduce_sd153;
  assign multm_reduce_ms154 = multm_reduce_add3b0_xor3b_wx154 ^ multm_reduce_sd154;
  assign multm_reduce_ms155 = multm_reduce_add3b0_xor3b_wx155 ^ multm_reduce_sd155;
  assign multm_reduce_ms156 = multm_reduce_add3b0_xor3b_wx156 ^ multm_reduce_sd156;
  assign multm_reduce_ms157 = multm_reduce_add3b0_xor3b_wx157 ^ multm_reduce_sd157;
  assign multm_reduce_ms158 = multm_reduce_add3b0_xor3b_wx158 ^ multm_reduce_sd158;
  assign multm_reduce_ms159 = multm_reduce_add3b0_xor3b_wx159 ^ multm_reduce_sd159;
  assign multm_reduce_ms160 = multm_reduce_add3b0_xor3b_wx160 ^ multm_reduce_sd160;
  assign multm_reduce_ms161 = multm_reduce_add3b0_xor3b_wx161 ^ multm_reduce_sd161;
  assign multm_reduce_ms162 = multm_reduce_add3b0_xor3b_wx162 ^ multm_reduce_sd162;
  assign multm_reduce_ms163 = multm_reduce_add3b0_xor3b_wx163 ^ multm_reduce_sd163;
  assign multm_reduce_ms164 = multm_reduce_add3b0_xor3b_wx164 ^ multm_reduce_sd164;
  assign multm_reduce_ms165 = multm_reduce_add3b0_xor3b_wx165 ^ multm_reduce_sd165;
  assign multm_reduce_ms166 = multm_reduce_add3b0_xor3b_wx166 ^ multm_reduce_sd166;
  assign multm_reduce_ms167 = multm_reduce_add3b0_xor3b_wx167 ^ multm_reduce_sd167;
  assign multm_reduce_ms168 = multm_reduce_add3b0_xor3b_wx168 ^ multm_reduce_sd168;
  assign multm_reduce_ms169 = multm_reduce_add3b0_xor3b_wx169 ^ multm_reduce_sd169;
  assign multm_reduce_ms170 = multm_reduce_add3b0_xor3b_wx170 ^ multm_reduce_sd170;
  assign multm_reduce_ms171 = multm_reduce_add3b0_xor3b_wx171 ^ multm_reduce_sd171;
  assign multm_reduce_ms172 = multm_reduce_add3b0_xor3b_wx172 ^ multm_reduce_sd172;
  assign multm_reduce_ms173 = multm_reduce_add3b0_xor3b_wx173 ^ multm_reduce_sd173;
  assign multm_reduce_ms174 = multm_reduce_add3b0_xor3b_wx174 ^ multm_reduce_sd174;
  assign multm_reduce_ms175 = multm_reduce_add3b0_xor3b_wx175 ^ multm_reduce_sd175;
  assign multm_reduce_ms176 = multm_reduce_add3b0_xor3b_wx176 ^ multm_reduce_sd176;
  assign multm_reduce_ms177 = multm_reduce_add3b0_xor3b_wx177 ^ multm_reduce_sd177;
  assign multm_reduce_ms178 = multm_reduce_add3b0_xor3b_wx178 ^ multm_reduce_sd178;
  assign multm_reduce_ms179 = multm_reduce_add3b0_xor3b_wx179 ^ multm_reduce_sd179;
  assign multm_reduce_ms180 = multm_reduce_add3b0_xor3b_wx180 ^ multm_reduce_sd180;
  assign multm_reduce_ms181 = multm_reduce_add3b0_xor3b_wx181 ^ multm_reduce_sd181;
  assign multm_reduce_ms182 = multm_reduce_add3b0_xor3b_wx182 ^ multm_reduce_sd182;
  assign multm_reduce_ms183 = multm_reduce_sa183 ^ multm_reduce_sd183;
  assign multm_reduce_mulb0_add3_maj3_or3_wx = multm_reduce_mulb0_add3_maj3_wx | multm_reduce_mulb0_add3_maj3_wy;
  assign multm_reduce_mulb0_add3_maj3_wx = multm_reduce_sa5 & multm_reduce_mulb0_cq184;
  assign multm_reduce_mulb0_add3_maj3_wy = multm_reduce_sa5 & multm_reduce_mulb0_pc184;
  assign multm_reduce_mulb0_add3_maj3_xy = multm_reduce_mulb0_cq184 & multm_reduce_mulb0_pc184;
  assign multm_reduce_mulb0_add3_xor3_wx = multm_reduce_sa5 ^ multm_reduce_mulb0_cq184;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx2 = multm_reduce_mulb0_add3b_maj3b_wx2 | multm_reduce_mulb0_add3b_maj3b_wy2;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx4 = multm_reduce_mulb0_add3b_maj3b_wx4 | multm_reduce_mulb0_add3b_maj3b_wy4;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx8 = multm_reduce_mulb0_add3b_maj3b_wx8 | multm_reduce_mulb0_add3b_maj3b_wy8;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx9 = multm_reduce_mulb0_add3b_maj3b_wx9 | multm_reduce_mulb0_add3b_maj3b_wy9;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx12 = multm_reduce_mulb0_add3b_maj3b_wx12 | multm_reduce_mulb0_add3b_maj3b_wy12;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx15 = multm_reduce_mulb0_add3b_maj3b_wx15 | multm_reduce_mulb0_add3b_maj3b_wy15;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx16 = multm_reduce_mulb0_add3b_maj3b_wx16 | multm_reduce_mulb0_add3b_maj3b_wy16;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx17 = multm_reduce_mulb0_add3b_maj3b_wx17 | multm_reduce_mulb0_add3b_maj3b_wy17;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx18 = multm_reduce_mulb0_add3b_maj3b_wx18 | multm_reduce_mulb0_add3b_maj3b_wy18;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx19 = multm_reduce_mulb0_add3b_maj3b_wx19 | multm_reduce_mulb0_add3b_maj3b_wy19;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx20 = multm_reduce_mulb0_add3b_maj3b_wx20 | multm_reduce_mulb0_add3b_maj3b_wy20;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx25 = multm_reduce_mulb0_add3b_maj3b_wx25 | multm_reduce_mulb0_add3b_maj3b_wy25;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx26 = multm_reduce_mulb0_add3b_maj3b_wx26 | multm_reduce_mulb0_add3b_maj3b_wy26;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx27 = multm_reduce_mulb0_add3b_maj3b_wx27 | multm_reduce_mulb0_add3b_maj3b_wy27;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx29 = multm_reduce_mulb0_add3b_maj3b_wx29 | multm_reduce_mulb0_add3b_maj3b_wy29;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx30 = multm_reduce_mulb0_add3b_maj3b_wx30 | multm_reduce_mulb0_add3b_maj3b_wy30;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx33 = multm_reduce_mulb0_add3b_maj3b_wx33 | multm_reduce_mulb0_add3b_maj3b_wy33;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx37 = multm_reduce_mulb0_add3b_maj3b_wx37 | multm_reduce_mulb0_add3b_maj3b_wy37;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx40 = multm_reduce_mulb0_add3b_maj3b_wx40 | multm_reduce_mulb0_add3b_maj3b_wy40;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx42 = multm_reduce_mulb0_add3b_maj3b_wx42 | multm_reduce_mulb0_add3b_maj3b_wy42;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx44 = multm_reduce_mulb0_add3b_maj3b_wx44 | multm_reduce_mulb0_add3b_maj3b_wy44;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx45 = multm_reduce_mulb0_add3b_maj3b_wx45 | multm_reduce_mulb0_add3b_maj3b_wy45;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx46 = multm_reduce_mulb0_add3b_maj3b_wx46 | multm_reduce_mulb0_add3b_maj3b_wy46;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx48 = multm_reduce_mulb0_add3b_maj3b_wx48 | multm_reduce_mulb0_add3b_maj3b_wy48;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx50 = multm_reduce_mulb0_add3b_maj3b_wx50 | multm_reduce_mulb0_add3b_maj3b_wy50;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx51 = multm_reduce_mulb0_add3b_maj3b_wx51 | multm_reduce_mulb0_add3b_maj3b_wy51;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx52 = multm_reduce_mulb0_add3b_maj3b_wx52 | multm_reduce_mulb0_add3b_maj3b_wy52;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx53 = multm_reduce_mulb0_add3b_maj3b_wx53 | multm_reduce_mulb0_add3b_maj3b_wy53;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx54 = multm_reduce_mulb0_add3b_maj3b_wx54 | multm_reduce_mulb0_add3b_maj3b_wy54;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx56 = multm_reduce_mulb0_add3b_maj3b_wx56 | multm_reduce_mulb0_add3b_maj3b_wy56;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx57 = multm_reduce_mulb0_add3b_maj3b_wx57 | multm_reduce_mulb0_add3b_maj3b_wy57;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx58 = multm_reduce_mulb0_add3b_maj3b_wx58 | multm_reduce_mulb0_add3b_maj3b_wy58;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx60 = multm_reduce_mulb0_add3b_maj3b_wx60 | multm_reduce_mulb0_add3b_maj3b_wy60;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx61 = multm_reduce_mulb0_add3b_maj3b_wx61 | multm_reduce_mulb0_add3b_maj3b_wy61;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx62 = multm_reduce_mulb0_add3b_maj3b_wx62 | multm_reduce_mulb0_add3b_maj3b_wy62;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx63 = multm_reduce_mulb0_add3b_maj3b_wx63 | multm_reduce_mulb0_add3b_maj3b_wy63;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx65 = multm_reduce_mulb0_add3b_maj3b_wx65 | multm_reduce_mulb0_add3b_maj3b_wy65;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx66 = multm_reduce_mulb0_add3b_maj3b_wx66 | multm_reduce_mulb0_add3b_maj3b_wy66;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx67 = multm_reduce_mulb0_add3b_maj3b_wx67 | multm_reduce_mulb0_add3b_maj3b_wy67;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx69 = multm_reduce_mulb0_add3b_maj3b_wx69 | multm_reduce_mulb0_add3b_maj3b_wy69;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx72 = multm_reduce_mulb0_add3b_maj3b_wx72 | multm_reduce_mulb0_add3b_maj3b_wy72;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx73 = multm_reduce_mulb0_add3b_maj3b_wx73 | multm_reduce_mulb0_add3b_maj3b_wy73;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx76 = multm_reduce_mulb0_add3b_maj3b_wx76 | multm_reduce_mulb0_add3b_maj3b_wy76;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx78 = multm_reduce_mulb0_add3b_maj3b_wx78 | multm_reduce_mulb0_add3b_maj3b_wy78;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx80 = multm_reduce_mulb0_add3b_maj3b_wx80 | multm_reduce_mulb0_add3b_maj3b_wy80;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx82 = multm_reduce_mulb0_add3b_maj3b_wx82 | multm_reduce_mulb0_add3b_maj3b_wy82;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx83 = multm_reduce_mulb0_add3b_maj3b_wx83 | multm_reduce_mulb0_add3b_maj3b_wy83;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx84 = multm_reduce_mulb0_add3b_maj3b_wx84 | multm_reduce_mulb0_add3b_maj3b_wy84;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx87 = multm_reduce_mulb0_add3b_maj3b_wx87 | multm_reduce_mulb0_add3b_maj3b_wy87;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx91 = multm_reduce_mulb0_add3b_maj3b_wx91 | multm_reduce_mulb0_add3b_maj3b_wy91;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx92 = multm_reduce_mulb0_add3b_maj3b_wx92 | multm_reduce_mulb0_add3b_maj3b_wy92;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx95 = multm_reduce_mulb0_add3b_maj3b_wx95 | multm_reduce_mulb0_add3b_maj3b_wy95;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx102 = multm_reduce_mulb0_add3b_maj3b_wx102 | multm_reduce_mulb0_add3b_maj3b_wy102;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx103 = multm_reduce_mulb0_add3b_maj3b_wx103 | multm_reduce_mulb0_add3b_maj3b_wy103;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx105 = multm_reduce_mulb0_add3b_maj3b_wx105 | multm_reduce_mulb0_add3b_maj3b_wy105;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx109 = multm_reduce_mulb0_add3b_maj3b_wx109 | multm_reduce_mulb0_add3b_maj3b_wy109;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx110 = multm_reduce_mulb0_add3b_maj3b_wx110 | multm_reduce_mulb0_add3b_maj3b_wy110;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx114 = multm_reduce_mulb0_add3b_maj3b_wx114 | multm_reduce_mulb0_add3b_maj3b_wy114;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx117 = multm_reduce_mulb0_add3b_maj3b_wx117 | multm_reduce_mulb0_add3b_maj3b_wy117;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx118 = multm_reduce_mulb0_add3b_maj3b_wx118 | multm_reduce_mulb0_add3b_maj3b_wy118;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx120 = multm_reduce_mulb0_add3b_maj3b_wx120 | multm_reduce_mulb0_add3b_maj3b_wy120;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx122 = multm_reduce_mulb0_add3b_maj3b_wx122 | multm_reduce_mulb0_add3b_maj3b_wy122;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx123 = multm_reduce_mulb0_add3b_maj3b_wx123 | multm_reduce_mulb0_add3b_maj3b_wy123;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx127 = multm_reduce_mulb0_add3b_maj3b_wx127 | multm_reduce_mulb0_add3b_maj3b_wy127;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx128 = multm_reduce_mulb0_add3b_maj3b_wx128 | multm_reduce_mulb0_add3b_maj3b_wy128;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx131 = multm_reduce_mulb0_add3b_maj3b_wx131 | multm_reduce_mulb0_add3b_maj3b_wy131;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx134 = multm_reduce_mulb0_add3b_maj3b_wx134 | multm_reduce_mulb0_add3b_maj3b_wy134;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx135 = multm_reduce_mulb0_add3b_maj3b_wx135 | multm_reduce_mulb0_add3b_maj3b_wy135;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx136 = multm_reduce_mulb0_add3b_maj3b_wx136 | multm_reduce_mulb0_add3b_maj3b_wy136;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx138 = multm_reduce_mulb0_add3b_maj3b_wx138 | multm_reduce_mulb0_add3b_maj3b_wy138;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx140 = multm_reduce_mulb0_add3b_maj3b_wx140 | multm_reduce_mulb0_add3b_maj3b_wy140;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx146 = multm_reduce_mulb0_add3b_maj3b_wx146 | multm_reduce_mulb0_add3b_maj3b_wy146;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx147 = multm_reduce_mulb0_add3b_maj3b_wx147 | multm_reduce_mulb0_add3b_maj3b_wy147;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx148 = multm_reduce_mulb0_add3b_maj3b_wx148 | multm_reduce_mulb0_add3b_maj3b_wy148;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx149 = multm_reduce_mulb0_add3b_maj3b_wx149 | multm_reduce_mulb0_add3b_maj3b_wy149;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx152 = multm_reduce_mulb0_add3b_maj3b_wx152 | multm_reduce_mulb0_add3b_maj3b_wy152;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx153 = multm_reduce_mulb0_add3b_maj3b_wx153 | multm_reduce_mulb0_add3b_maj3b_wy153;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx156 = multm_reduce_mulb0_add3b_maj3b_wx156 | multm_reduce_mulb0_add3b_maj3b_wy156;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx157 = multm_reduce_mulb0_add3b_maj3b_wx157 | multm_reduce_mulb0_add3b_maj3b_wy157;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx158 = multm_reduce_mulb0_add3b_maj3b_wx158 | multm_reduce_mulb0_add3b_maj3b_wy158;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx159 = multm_reduce_mulb0_add3b_maj3b_wx159 | multm_reduce_mulb0_add3b_maj3b_wy159;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx160 = multm_reduce_mulb0_add3b_maj3b_wx160 | multm_reduce_mulb0_add3b_maj3b_wy160;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx162 = multm_reduce_mulb0_add3b_maj3b_wx162 | multm_reduce_mulb0_add3b_maj3b_wy162;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx163 = multm_reduce_mulb0_add3b_maj3b_wx163 | multm_reduce_mulb0_add3b_maj3b_wy163;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx168 = multm_reduce_mulb0_add3b_maj3b_wx168 | multm_reduce_mulb0_add3b_maj3b_wy168;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx170 = multm_reduce_mulb0_add3b_maj3b_wx170 | multm_reduce_mulb0_add3b_maj3b_wy170;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx171 = multm_reduce_mulb0_add3b_maj3b_wx171 | multm_reduce_mulb0_add3b_maj3b_wy171;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx172 = multm_reduce_mulb0_add3b_maj3b_wx172 | multm_reduce_mulb0_add3b_maj3b_wy172;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx173 = multm_reduce_mulb0_add3b_maj3b_wx173 | multm_reduce_mulb0_add3b_maj3b_wy173;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx175 = multm_reduce_mulb0_add3b_maj3b_wx175 | multm_reduce_mulb0_add3b_maj3b_wy175;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx177 = multm_reduce_mulb0_add3b_maj3b_wx177 | multm_reduce_mulb0_add3b_maj3b_wy177;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx178 = multm_reduce_mulb0_add3b_maj3b_wx178 | multm_reduce_mulb0_add3b_maj3b_wy178;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx181 = multm_reduce_mulb0_add3b_maj3b_wx181 | multm_reduce_mulb0_add3b_maj3b_wy181;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx182 = multm_reduce_mulb0_add3b_maj3b_wx182 | multm_reduce_mulb0_add3b_maj3b_wy182;
  assign multm_reduce_mulb0_add3b_maj3b_or3b_wx183 = multm_reduce_mulb0_add3b_maj3b_wx183 | multm_reduce_mulb0_add3b_maj3b_wy183;
  assign multm_reduce_mulb0_add3b_maj3b_wx2 = multm_reduce_mulb0_sq3 & multm_reduce_mulb0_cq2;
  assign multm_reduce_mulb0_add3b_maj3b_wx4 = multm_reduce_mulb0_sq5 & multm_reduce_mulb0_cq4;
  assign multm_reduce_mulb0_add3b_maj3b_wx8 = multm_reduce_mulb0_sq9 & multm_reduce_mulb0_cq8;
  assign multm_reduce_mulb0_add3b_maj3b_wx9 = multm_reduce_mulb0_sq10 & multm_reduce_mulb0_cq9;
  assign multm_reduce_mulb0_add3b_maj3b_wx12 = multm_reduce_mulb0_sq13 & multm_reduce_mulb0_cq12;
  assign multm_reduce_mulb0_add3b_maj3b_wx15 = multm_reduce_mulb0_sq16 & multm_reduce_mulb0_cq15;
  assign multm_reduce_mulb0_add3b_maj3b_wx16 = multm_reduce_mulb0_sq17 & multm_reduce_mulb0_cq16;
  assign multm_reduce_mulb0_add3b_maj3b_wx17 = multm_reduce_mulb0_sq18 & multm_reduce_mulb0_cq17;
  assign multm_reduce_mulb0_add3b_maj3b_wx18 = multm_reduce_mulb0_sq19 & multm_reduce_mulb0_cq18;
  assign multm_reduce_mulb0_add3b_maj3b_wx19 = multm_reduce_mulb0_sq20 & multm_reduce_mulb0_cq19;
  assign multm_reduce_mulb0_add3b_maj3b_wx20 = multm_reduce_mulb0_sq21 & multm_reduce_mulb0_cq20;
  assign multm_reduce_mulb0_add3b_maj3b_wx25 = multm_reduce_mulb0_sq26 & multm_reduce_mulb0_cq25;
  assign multm_reduce_mulb0_add3b_maj3b_wx26 = multm_reduce_mulb0_sq27 & multm_reduce_mulb0_cq26;
  assign multm_reduce_mulb0_add3b_maj3b_wx27 = multm_reduce_mulb0_sq28 & multm_reduce_mulb0_cq27;
  assign multm_reduce_mulb0_add3b_maj3b_wx29 = multm_reduce_mulb0_sq30 & multm_reduce_mulb0_cq29;
  assign multm_reduce_mulb0_add3b_maj3b_wx30 = multm_reduce_mulb0_sq31 & multm_reduce_mulb0_cq30;
  assign multm_reduce_mulb0_add3b_maj3b_wx33 = multm_reduce_mulb0_sq34 & multm_reduce_mulb0_cq33;
  assign multm_reduce_mulb0_add3b_maj3b_wx37 = multm_reduce_mulb0_sq38 & multm_reduce_mulb0_cq37;
  assign multm_reduce_mulb0_add3b_maj3b_wx40 = multm_reduce_mulb0_sq41 & multm_reduce_mulb0_cq40;
  assign multm_reduce_mulb0_add3b_maj3b_wx42 = multm_reduce_mulb0_sq43 & multm_reduce_mulb0_cq42;
  assign multm_reduce_mulb0_add3b_maj3b_wx44 = multm_reduce_mulb0_sq45 & multm_reduce_mulb0_cq44;
  assign multm_reduce_mulb0_add3b_maj3b_wx45 = multm_reduce_mulb0_sq46 & multm_reduce_mulb0_cq45;
  assign multm_reduce_mulb0_add3b_maj3b_wx46 = multm_reduce_mulb0_sq47 & multm_reduce_mulb0_cq46;
  assign multm_reduce_mulb0_add3b_maj3b_wx48 = multm_reduce_mulb0_sq49 & multm_reduce_mulb0_cq48;
  assign multm_reduce_mulb0_add3b_maj3b_wx50 = multm_reduce_mulb0_sq51 & multm_reduce_mulb0_cq50;
  assign multm_reduce_mulb0_add3b_maj3b_wx51 = multm_reduce_mulb0_sq52 & multm_reduce_mulb0_cq51;
  assign multm_reduce_mulb0_add3b_maj3b_wx52 = multm_reduce_mulb0_sq53 & multm_reduce_mulb0_cq52;
  assign multm_reduce_mulb0_add3b_maj3b_wx53 = multm_reduce_mulb0_sq54 & multm_reduce_mulb0_cq53;
  assign multm_reduce_mulb0_add3b_maj3b_wx54 = multm_reduce_mulb0_sq55 & multm_reduce_mulb0_cq54;
  assign multm_reduce_mulb0_add3b_maj3b_wx56 = multm_reduce_mulb0_sq57 & multm_reduce_mulb0_cq56;
  assign multm_reduce_mulb0_add3b_maj3b_wx57 = multm_reduce_mulb0_sq58 & multm_reduce_mulb0_cq57;
  assign multm_reduce_mulb0_add3b_maj3b_wx58 = multm_reduce_mulb0_sq59 & multm_reduce_mulb0_cq58;
  assign multm_reduce_mulb0_add3b_maj3b_wx60 = multm_reduce_mulb0_sq61 & multm_reduce_mulb0_cq60;
  assign multm_reduce_mulb0_add3b_maj3b_wx61 = multm_reduce_mulb0_sq62 & multm_reduce_mulb0_cq61;
  assign multm_reduce_mulb0_add3b_maj3b_wx62 = multm_reduce_mulb0_sq63 & multm_reduce_mulb0_cq62;
  assign multm_reduce_mulb0_add3b_maj3b_wx63 = multm_reduce_mulb0_sq64 & multm_reduce_mulb0_cq63;
  assign multm_reduce_mulb0_add3b_maj3b_wx65 = multm_reduce_mulb0_sq66 & multm_reduce_mulb0_cq65;
  assign multm_reduce_mulb0_add3b_maj3b_wx66 = multm_reduce_mulb0_sq67 & multm_reduce_mulb0_cq66;
  assign multm_reduce_mulb0_add3b_maj3b_wx67 = multm_reduce_mulb0_sq68 & multm_reduce_mulb0_cq67;
  assign multm_reduce_mulb0_add3b_maj3b_wx69 = multm_reduce_mulb0_sq70 & multm_reduce_mulb0_cq69;
  assign multm_reduce_mulb0_add3b_maj3b_wx72 = multm_reduce_mulb0_sq73 & multm_reduce_mulb0_cq72;
  assign multm_reduce_mulb0_add3b_maj3b_wx73 = multm_reduce_mulb0_sq74 & multm_reduce_mulb0_cq73;
  assign multm_reduce_mulb0_add3b_maj3b_wx76 = multm_reduce_mulb0_sq77 & multm_reduce_mulb0_cq76;
  assign multm_reduce_mulb0_add3b_maj3b_wx78 = multm_reduce_mulb0_sq79 & multm_reduce_mulb0_cq78;
  assign multm_reduce_mulb0_add3b_maj3b_wx80 = multm_reduce_mulb0_sq81 & multm_reduce_mulb0_cq80;
  assign multm_reduce_mulb0_add3b_maj3b_wx82 = multm_reduce_mulb0_sq83 & multm_reduce_mulb0_cq82;
  assign multm_reduce_mulb0_add3b_maj3b_wx83 = multm_reduce_mulb0_sq84 & multm_reduce_mulb0_cq83;
  assign multm_reduce_mulb0_add3b_maj3b_wx84 = multm_reduce_mulb0_sq85 & multm_reduce_mulb0_cq84;
  assign multm_reduce_mulb0_add3b_maj3b_wx87 = multm_reduce_mulb0_sq88 & multm_reduce_mulb0_cq87;
  assign multm_reduce_mulb0_add3b_maj3b_wx91 = multm_reduce_mulb0_sq92 & multm_reduce_mulb0_cq91;
  assign multm_reduce_mulb0_add3b_maj3b_wx92 = multm_reduce_mulb0_sq93 & multm_reduce_mulb0_cq92;
  assign multm_reduce_mulb0_add3b_maj3b_wx95 = multm_reduce_mulb0_sq96 & multm_reduce_mulb0_cq95;
  assign multm_reduce_mulb0_add3b_maj3b_wx102 = multm_reduce_mulb0_sq103 & multm_reduce_mulb0_cq102;
  assign multm_reduce_mulb0_add3b_maj3b_wx103 = multm_reduce_mulb0_sq104 & multm_reduce_mulb0_cq103;
  assign multm_reduce_mulb0_add3b_maj3b_wx105 = multm_reduce_mulb0_sq106 & multm_reduce_mulb0_cq105;
  assign multm_reduce_mulb0_add3b_maj3b_wx109 = multm_reduce_mulb0_sq110 & multm_reduce_mulb0_cq109;
  assign multm_reduce_mulb0_add3b_maj3b_wx110 = multm_reduce_mulb0_sq111 & multm_reduce_mulb0_cq110;
  assign multm_reduce_mulb0_add3b_maj3b_wx114 = multm_reduce_mulb0_sq115 & multm_reduce_mulb0_cq114;
  assign multm_reduce_mulb0_add3b_maj3b_wx117 = multm_reduce_mulb0_sq118 & multm_reduce_mulb0_cq117;
  assign multm_reduce_mulb0_add3b_maj3b_wx118 = multm_reduce_mulb0_sq119 & multm_reduce_mulb0_cq118;
  assign multm_reduce_mulb0_add3b_maj3b_wx120 = multm_reduce_mulb0_sq121 & multm_reduce_mulb0_cq120;
  assign multm_reduce_mulb0_add3b_maj3b_wx122 = multm_reduce_mulb0_sq123 & multm_reduce_mulb0_cq122;
  assign multm_reduce_mulb0_add3b_maj3b_wx123 = multm_reduce_mulb0_sq124 & multm_reduce_mulb0_cq123;
  assign multm_reduce_mulb0_add3b_maj3b_wx127 = multm_reduce_mulb0_sq128 & multm_reduce_mulb0_cq127;
  assign multm_reduce_mulb0_add3b_maj3b_wx128 = multm_reduce_mulb0_sq129 & multm_reduce_mulb0_cq128;
  assign multm_reduce_mulb0_add3b_maj3b_wx131 = multm_reduce_mulb0_sq132 & multm_reduce_mulb0_cq131;
  assign multm_reduce_mulb0_add3b_maj3b_wx134 = multm_reduce_mulb0_sq135 & multm_reduce_mulb0_cq134;
  assign multm_reduce_mulb0_add3b_maj3b_wx135 = multm_reduce_mulb0_sq136 & multm_reduce_mulb0_cq135;
  assign multm_reduce_mulb0_add3b_maj3b_wx136 = multm_reduce_mulb0_sq137 & multm_reduce_mulb0_cq136;
  assign multm_reduce_mulb0_add3b_maj3b_wx138 = multm_reduce_mulb0_sq139 & multm_reduce_mulb0_cq138;
  assign multm_reduce_mulb0_add3b_maj3b_wx140 = multm_reduce_mulb0_sq141 & multm_reduce_mulb0_cq140;
  assign multm_reduce_mulb0_add3b_maj3b_wx146 = multm_reduce_mulb0_sq147 & multm_reduce_mulb0_cq146;
  assign multm_reduce_mulb0_add3b_maj3b_wx147 = multm_reduce_mulb0_sq148 & multm_reduce_mulb0_cq147;
  assign multm_reduce_mulb0_add3b_maj3b_wx148 = multm_reduce_mulb0_sq149 & multm_reduce_mulb0_cq148;
  assign multm_reduce_mulb0_add3b_maj3b_wx149 = multm_reduce_mulb0_sq150 & multm_reduce_mulb0_cq149;
  assign multm_reduce_mulb0_add3b_maj3b_wx152 = multm_reduce_mulb0_sq153 & multm_reduce_mulb0_cq152;
  assign multm_reduce_mulb0_add3b_maj3b_wx153 = multm_reduce_mulb0_sq154 & multm_reduce_mulb0_cq153;
  assign multm_reduce_mulb0_add3b_maj3b_wx156 = multm_reduce_mulb0_sq157 & multm_reduce_mulb0_cq156;
  assign multm_reduce_mulb0_add3b_maj3b_wx157 = multm_reduce_mulb0_sq158 & multm_reduce_mulb0_cq157;
  assign multm_reduce_mulb0_add3b_maj3b_wx158 = multm_reduce_mulb0_sq159 & multm_reduce_mulb0_cq158;
  assign multm_reduce_mulb0_add3b_maj3b_wx159 = multm_reduce_mulb0_sq160 & multm_reduce_mulb0_cq159;
  assign multm_reduce_mulb0_add3b_maj3b_wx160 = multm_reduce_mulb0_sq161 & multm_reduce_mulb0_cq160;
  assign multm_reduce_mulb0_add3b_maj3b_wx162 = multm_reduce_mulb0_sq163 & multm_reduce_mulb0_cq162;
  assign multm_reduce_mulb0_add3b_maj3b_wx163 = multm_reduce_mulb0_sq164 & multm_reduce_mulb0_cq163;
  assign multm_reduce_mulb0_add3b_maj3b_wx168 = multm_reduce_mulb0_sq169 & multm_reduce_mulb0_cq168;
  assign multm_reduce_mulb0_add3b_maj3b_wx170 = multm_reduce_mulb0_sq171 & multm_reduce_mulb0_cq170;
  assign multm_reduce_mulb0_add3b_maj3b_wx171 = multm_reduce_mulb0_sq172 & multm_reduce_mulb0_cq171;
  assign multm_reduce_mulb0_add3b_maj3b_wx172 = multm_reduce_mulb0_sq173 & multm_reduce_mulb0_cq172;
  assign multm_reduce_mulb0_add3b_maj3b_wx173 = multm_reduce_mulb0_sq174 & multm_reduce_mulb0_cq173;
  assign multm_reduce_mulb0_add3b_maj3b_wx175 = multm_reduce_mulb0_sq176 & multm_reduce_mulb0_cq175;
  assign multm_reduce_mulb0_add3b_maj3b_wx177 = multm_reduce_mulb0_sq178 & multm_reduce_mulb0_cq177;
  assign multm_reduce_mulb0_add3b_maj3b_wx178 = multm_reduce_mulb0_sq179 & multm_reduce_mulb0_cq178;
  assign multm_reduce_mulb0_add3b_maj3b_wx181 = multm_reduce_mulb0_sq182 & multm_reduce_mulb0_cq181;
  assign multm_reduce_mulb0_add3b_maj3b_wx182 = multm_reduce_mulb0_sq183 & multm_reduce_mulb0_cq182;
  assign multm_reduce_mulb0_add3b_maj3b_wx183 = multm_reduce_mulb0_sq184 & multm_reduce_mulb0_cq183;
  assign multm_reduce_mulb0_add3b_maj3b_wy2 = multm_reduce_mulb0_sq3 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy4 = multm_reduce_mulb0_sq5 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy8 = multm_reduce_mulb0_sq9 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy9 = multm_reduce_mulb0_sq10 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy12 = multm_reduce_mulb0_sq13 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy15 = multm_reduce_mulb0_sq16 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy16 = multm_reduce_mulb0_sq17 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy17 = multm_reduce_mulb0_sq18 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy18 = multm_reduce_mulb0_sq19 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy19 = multm_reduce_mulb0_sq20 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy20 = multm_reduce_mulb0_sq21 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy25 = multm_reduce_mulb0_sq26 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy26 = multm_reduce_mulb0_sq27 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy27 = multm_reduce_mulb0_sq28 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy29 = multm_reduce_mulb0_sq30 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy30 = multm_reduce_mulb0_sq31 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy33 = multm_reduce_mulb0_sq34 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy37 = multm_reduce_mulb0_sq38 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy40 = multm_reduce_mulb0_sq41 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy42 = multm_reduce_mulb0_sq43 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy44 = multm_reduce_mulb0_sq45 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy45 = multm_reduce_mulb0_sq46 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy46 = multm_reduce_mulb0_sq47 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy48 = multm_reduce_mulb0_sq49 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy50 = multm_reduce_mulb0_sq51 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy51 = multm_reduce_mulb0_sq52 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy52 = multm_reduce_mulb0_sq53 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy53 = multm_reduce_mulb0_sq54 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy54 = multm_reduce_mulb0_sq55 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy56 = multm_reduce_mulb0_sq57 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy57 = multm_reduce_mulb0_sq58 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy58 = multm_reduce_mulb0_sq59 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy60 = multm_reduce_mulb0_sq61 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy61 = multm_reduce_mulb0_sq62 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy62 = multm_reduce_mulb0_sq63 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy63 = multm_reduce_mulb0_sq64 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy65 = multm_reduce_mulb0_sq66 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy66 = multm_reduce_mulb0_sq67 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy67 = multm_reduce_mulb0_sq68 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy69 = multm_reduce_mulb0_sq70 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy72 = multm_reduce_mulb0_sq73 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy73 = multm_reduce_mulb0_sq74 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy76 = multm_reduce_mulb0_sq77 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy78 = multm_reduce_mulb0_sq79 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy80 = multm_reduce_mulb0_sq81 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy82 = multm_reduce_mulb0_sq83 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy83 = multm_reduce_mulb0_sq84 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy84 = multm_reduce_mulb0_sq85 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy87 = multm_reduce_mulb0_sq88 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy91 = multm_reduce_mulb0_sq92 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy92 = multm_reduce_mulb0_sq93 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy95 = multm_reduce_mulb0_sq96 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy102 = multm_reduce_mulb0_sq103 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy103 = multm_reduce_mulb0_sq104 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy105 = multm_reduce_mulb0_sq106 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy109 = multm_reduce_mulb0_sq110 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy110 = multm_reduce_mulb0_sq111 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy114 = multm_reduce_mulb0_sq115 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy117 = multm_reduce_mulb0_sq118 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy118 = multm_reduce_mulb0_sq119 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy120 = multm_reduce_mulb0_sq121 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy122 = multm_reduce_mulb0_sq123 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy123 = multm_reduce_mulb0_sq124 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy127 = multm_reduce_mulb0_sq128 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy128 = multm_reduce_mulb0_sq129 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy131 = multm_reduce_mulb0_sq132 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy134 = multm_reduce_mulb0_sq135 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy135 = multm_reduce_mulb0_sq136 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy136 = multm_reduce_mulb0_sq137 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy138 = multm_reduce_mulb0_sq139 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy140 = multm_reduce_mulb0_sq141 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy146 = multm_reduce_mulb0_sq147 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy147 = multm_reduce_mulb0_sq148 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy148 = multm_reduce_mulb0_sq149 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy149 = multm_reduce_mulb0_sq150 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy152 = multm_reduce_mulb0_sq153 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy153 = multm_reduce_mulb0_sq154 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy156 = multm_reduce_mulb0_sq157 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy157 = multm_reduce_mulb0_sq158 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy158 = multm_reduce_mulb0_sq159 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy159 = multm_reduce_mulb0_sq160 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy160 = multm_reduce_mulb0_sq161 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy162 = multm_reduce_mulb0_sq163 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy163 = multm_reduce_mulb0_sq164 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy168 = multm_reduce_mulb0_sq169 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy170 = multm_reduce_mulb0_sq171 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy171 = multm_reduce_mulb0_sq172 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy172 = multm_reduce_mulb0_sq173 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy173 = multm_reduce_mulb0_sq174 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy175 = multm_reduce_mulb0_sq176 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy177 = multm_reduce_mulb0_sq178 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy178 = multm_reduce_mulb0_sq179 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy181 = multm_reduce_mulb0_sq182 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy182 = multm_reduce_mulb0_sq183 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_wy183 = multm_reduce_mulb0_sq184 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy2 = multm_reduce_mulb0_cq2 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy4 = multm_reduce_mulb0_cq4 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy8 = multm_reduce_mulb0_cq8 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy9 = multm_reduce_mulb0_cq9 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy12 = multm_reduce_mulb0_cq12 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy15 = multm_reduce_mulb0_cq15 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy16 = multm_reduce_mulb0_cq16 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy17 = multm_reduce_mulb0_cq17 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy18 = multm_reduce_mulb0_cq18 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy19 = multm_reduce_mulb0_cq19 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy20 = multm_reduce_mulb0_cq20 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy25 = multm_reduce_mulb0_cq25 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy26 = multm_reduce_mulb0_cq26 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy27 = multm_reduce_mulb0_cq27 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy29 = multm_reduce_mulb0_cq29 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy30 = multm_reduce_mulb0_cq30 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy33 = multm_reduce_mulb0_cq33 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy37 = multm_reduce_mulb0_cq37 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy40 = multm_reduce_mulb0_cq40 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy42 = multm_reduce_mulb0_cq42 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy44 = multm_reduce_mulb0_cq44 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy45 = multm_reduce_mulb0_cq45 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy46 = multm_reduce_mulb0_cq46 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy48 = multm_reduce_mulb0_cq48 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy50 = multm_reduce_mulb0_cq50 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy51 = multm_reduce_mulb0_cq51 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy52 = multm_reduce_mulb0_cq52 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy53 = multm_reduce_mulb0_cq53 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy54 = multm_reduce_mulb0_cq54 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy56 = multm_reduce_mulb0_cq56 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy57 = multm_reduce_mulb0_cq57 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy58 = multm_reduce_mulb0_cq58 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy60 = multm_reduce_mulb0_cq60 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy61 = multm_reduce_mulb0_cq61 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy62 = multm_reduce_mulb0_cq62 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy63 = multm_reduce_mulb0_cq63 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy65 = multm_reduce_mulb0_cq65 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy66 = multm_reduce_mulb0_cq66 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy67 = multm_reduce_mulb0_cq67 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy69 = multm_reduce_mulb0_cq69 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy72 = multm_reduce_mulb0_cq72 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy73 = multm_reduce_mulb0_cq73 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy76 = multm_reduce_mulb0_cq76 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy78 = multm_reduce_mulb0_cq78 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy80 = multm_reduce_mulb0_cq80 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy82 = multm_reduce_mulb0_cq82 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy83 = multm_reduce_mulb0_cq83 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy84 = multm_reduce_mulb0_cq84 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy87 = multm_reduce_mulb0_cq87 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy91 = multm_reduce_mulb0_cq91 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy92 = multm_reduce_mulb0_cq92 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy95 = multm_reduce_mulb0_cq95 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy102 = multm_reduce_mulb0_cq102 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy103 = multm_reduce_mulb0_cq103 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy105 = multm_reduce_mulb0_cq105 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy109 = multm_reduce_mulb0_cq109 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy110 = multm_reduce_mulb0_cq110 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy114 = multm_reduce_mulb0_cq114 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy117 = multm_reduce_mulb0_cq117 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy118 = multm_reduce_mulb0_cq118 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy120 = multm_reduce_mulb0_cq120 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy122 = multm_reduce_mulb0_cq122 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy123 = multm_reduce_mulb0_cq123 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy127 = multm_reduce_mulb0_cq127 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy128 = multm_reduce_mulb0_cq128 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy131 = multm_reduce_mulb0_cq131 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy134 = multm_reduce_mulb0_cq134 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy135 = multm_reduce_mulb0_cq135 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy136 = multm_reduce_mulb0_cq136 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy138 = multm_reduce_mulb0_cq138 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy140 = multm_reduce_mulb0_cq140 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy146 = multm_reduce_mulb0_cq146 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy147 = multm_reduce_mulb0_cq147 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy148 = multm_reduce_mulb0_cq148 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy149 = multm_reduce_mulb0_cq149 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy152 = multm_reduce_mulb0_cq152 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy153 = multm_reduce_mulb0_cq153 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy156 = multm_reduce_mulb0_cq156 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy157 = multm_reduce_mulb0_cq157 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy158 = multm_reduce_mulb0_cq158 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy159 = multm_reduce_mulb0_cq159 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy160 = multm_reduce_mulb0_cq160 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy162 = multm_reduce_mulb0_cq162 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy163 = multm_reduce_mulb0_cq163 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy168 = multm_reduce_mulb0_cq168 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy170 = multm_reduce_mulb0_cq170 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy171 = multm_reduce_mulb0_cq171 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy172 = multm_reduce_mulb0_cq172 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy173 = multm_reduce_mulb0_cq173 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy175 = multm_reduce_mulb0_cq175 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy177 = multm_reduce_mulb0_cq177 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy178 = multm_reduce_mulb0_cq178 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy181 = multm_reduce_mulb0_cq181 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy182 = multm_reduce_mulb0_cq182 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_maj3b_xy183 = multm_reduce_mulb0_cq183 & multm_reduce_sa5;
  assign multm_reduce_mulb0_add3b_xor3b_wx2 = multm_reduce_mulb0_sq3 ^ multm_reduce_mulb0_cq2;
  assign multm_reduce_mulb0_add3b_xor3b_wx4 = multm_reduce_mulb0_sq5 ^ multm_reduce_mulb0_cq4;
  assign multm_reduce_mulb0_add3b_xor3b_wx8 = multm_reduce_mulb0_sq9 ^ multm_reduce_mulb0_cq8;
  assign multm_reduce_mulb0_add3b_xor3b_wx9 = multm_reduce_mulb0_sq10 ^ multm_reduce_mulb0_cq9;
  assign multm_reduce_mulb0_add3b_xor3b_wx12 = multm_reduce_mulb0_sq13 ^ multm_reduce_mulb0_cq12;
  assign multm_reduce_mulb0_add3b_xor3b_wx15 = multm_reduce_mulb0_sq16 ^ multm_reduce_mulb0_cq15;
  assign multm_reduce_mulb0_add3b_xor3b_wx16 = multm_reduce_mulb0_sq17 ^ multm_reduce_mulb0_cq16;
  assign multm_reduce_mulb0_add3b_xor3b_wx17 = multm_reduce_mulb0_sq18 ^ multm_reduce_mulb0_cq17;
  assign multm_reduce_mulb0_add3b_xor3b_wx18 = multm_reduce_mulb0_sq19 ^ multm_reduce_mulb0_cq18;
  assign multm_reduce_mulb0_add3b_xor3b_wx19 = multm_reduce_mulb0_sq20 ^ multm_reduce_mulb0_cq19;
  assign multm_reduce_mulb0_add3b_xor3b_wx20 = multm_reduce_mulb0_sq21 ^ multm_reduce_mulb0_cq20;
  assign multm_reduce_mulb0_add3b_xor3b_wx25 = multm_reduce_mulb0_sq26 ^ multm_reduce_mulb0_cq25;
  assign multm_reduce_mulb0_add3b_xor3b_wx26 = multm_reduce_mulb0_sq27 ^ multm_reduce_mulb0_cq26;
  assign multm_reduce_mulb0_add3b_xor3b_wx27 = multm_reduce_mulb0_sq28 ^ multm_reduce_mulb0_cq27;
  assign multm_reduce_mulb0_add3b_xor3b_wx29 = multm_reduce_mulb0_sq30 ^ multm_reduce_mulb0_cq29;
  assign multm_reduce_mulb0_add3b_xor3b_wx30 = multm_reduce_mulb0_sq31 ^ multm_reduce_mulb0_cq30;
  assign multm_reduce_mulb0_add3b_xor3b_wx33 = multm_reduce_mulb0_sq34 ^ multm_reduce_mulb0_cq33;
  assign multm_reduce_mulb0_add3b_xor3b_wx37 = multm_reduce_mulb0_sq38 ^ multm_reduce_mulb0_cq37;
  assign multm_reduce_mulb0_add3b_xor3b_wx40 = multm_reduce_mulb0_sq41 ^ multm_reduce_mulb0_cq40;
  assign multm_reduce_mulb0_add3b_xor3b_wx42 = multm_reduce_mulb0_sq43 ^ multm_reduce_mulb0_cq42;
  assign multm_reduce_mulb0_add3b_xor3b_wx44 = multm_reduce_mulb0_sq45 ^ multm_reduce_mulb0_cq44;
  assign multm_reduce_mulb0_add3b_xor3b_wx45 = multm_reduce_mulb0_sq46 ^ multm_reduce_mulb0_cq45;
  assign multm_reduce_mulb0_add3b_xor3b_wx46 = multm_reduce_mulb0_sq47 ^ multm_reduce_mulb0_cq46;
  assign multm_reduce_mulb0_add3b_xor3b_wx48 = multm_reduce_mulb0_sq49 ^ multm_reduce_mulb0_cq48;
  assign multm_reduce_mulb0_add3b_xor3b_wx50 = multm_reduce_mulb0_sq51 ^ multm_reduce_mulb0_cq50;
  assign multm_reduce_mulb0_add3b_xor3b_wx51 = multm_reduce_mulb0_sq52 ^ multm_reduce_mulb0_cq51;
  assign multm_reduce_mulb0_add3b_xor3b_wx52 = multm_reduce_mulb0_sq53 ^ multm_reduce_mulb0_cq52;
  assign multm_reduce_mulb0_add3b_xor3b_wx53 = multm_reduce_mulb0_sq54 ^ multm_reduce_mulb0_cq53;
  assign multm_reduce_mulb0_add3b_xor3b_wx54 = multm_reduce_mulb0_sq55 ^ multm_reduce_mulb0_cq54;
  assign multm_reduce_mulb0_add3b_xor3b_wx56 = multm_reduce_mulb0_sq57 ^ multm_reduce_mulb0_cq56;
  assign multm_reduce_mulb0_add3b_xor3b_wx57 = multm_reduce_mulb0_sq58 ^ multm_reduce_mulb0_cq57;
  assign multm_reduce_mulb0_add3b_xor3b_wx58 = multm_reduce_mulb0_sq59 ^ multm_reduce_mulb0_cq58;
  assign multm_reduce_mulb0_add3b_xor3b_wx60 = multm_reduce_mulb0_sq61 ^ multm_reduce_mulb0_cq60;
  assign multm_reduce_mulb0_add3b_xor3b_wx61 = multm_reduce_mulb0_sq62 ^ multm_reduce_mulb0_cq61;
  assign multm_reduce_mulb0_add3b_xor3b_wx62 = multm_reduce_mulb0_sq63 ^ multm_reduce_mulb0_cq62;
  assign multm_reduce_mulb0_add3b_xor3b_wx63 = multm_reduce_mulb0_sq64 ^ multm_reduce_mulb0_cq63;
  assign multm_reduce_mulb0_add3b_xor3b_wx65 = multm_reduce_mulb0_sq66 ^ multm_reduce_mulb0_cq65;
  assign multm_reduce_mulb0_add3b_xor3b_wx66 = multm_reduce_mulb0_sq67 ^ multm_reduce_mulb0_cq66;
  assign multm_reduce_mulb0_add3b_xor3b_wx67 = multm_reduce_mulb0_sq68 ^ multm_reduce_mulb0_cq67;
  assign multm_reduce_mulb0_add3b_xor3b_wx69 = multm_reduce_mulb0_sq70 ^ multm_reduce_mulb0_cq69;
  assign multm_reduce_mulb0_add3b_xor3b_wx72 = multm_reduce_mulb0_sq73 ^ multm_reduce_mulb0_cq72;
  assign multm_reduce_mulb0_add3b_xor3b_wx73 = multm_reduce_mulb0_sq74 ^ multm_reduce_mulb0_cq73;
  assign multm_reduce_mulb0_add3b_xor3b_wx76 = multm_reduce_mulb0_sq77 ^ multm_reduce_mulb0_cq76;
  assign multm_reduce_mulb0_add3b_xor3b_wx78 = multm_reduce_mulb0_sq79 ^ multm_reduce_mulb0_cq78;
  assign multm_reduce_mulb0_add3b_xor3b_wx80 = multm_reduce_mulb0_sq81 ^ multm_reduce_mulb0_cq80;
  assign multm_reduce_mulb0_add3b_xor3b_wx82 = multm_reduce_mulb0_sq83 ^ multm_reduce_mulb0_cq82;
  assign multm_reduce_mulb0_add3b_xor3b_wx83 = multm_reduce_mulb0_sq84 ^ multm_reduce_mulb0_cq83;
  assign multm_reduce_mulb0_add3b_xor3b_wx84 = multm_reduce_mulb0_sq85 ^ multm_reduce_mulb0_cq84;
  assign multm_reduce_mulb0_add3b_xor3b_wx87 = multm_reduce_mulb0_sq88 ^ multm_reduce_mulb0_cq87;
  assign multm_reduce_mulb0_add3b_xor3b_wx91 = multm_reduce_mulb0_sq92 ^ multm_reduce_mulb0_cq91;
  assign multm_reduce_mulb0_add3b_xor3b_wx92 = multm_reduce_mulb0_sq93 ^ multm_reduce_mulb0_cq92;
  assign multm_reduce_mulb0_add3b_xor3b_wx95 = multm_reduce_mulb0_sq96 ^ multm_reduce_mulb0_cq95;
  assign multm_reduce_mulb0_add3b_xor3b_wx102 = multm_reduce_mulb0_sq103 ^ multm_reduce_mulb0_cq102;
  assign multm_reduce_mulb0_add3b_xor3b_wx103 = multm_reduce_mulb0_sq104 ^ multm_reduce_mulb0_cq103;
  assign multm_reduce_mulb0_add3b_xor3b_wx105 = multm_reduce_mulb0_sq106 ^ multm_reduce_mulb0_cq105;
  assign multm_reduce_mulb0_add3b_xor3b_wx109 = multm_reduce_mulb0_sq110 ^ multm_reduce_mulb0_cq109;
  assign multm_reduce_mulb0_add3b_xor3b_wx110 = multm_reduce_mulb0_sq111 ^ multm_reduce_mulb0_cq110;
  assign multm_reduce_mulb0_add3b_xor3b_wx114 = multm_reduce_mulb0_sq115 ^ multm_reduce_mulb0_cq114;
  assign multm_reduce_mulb0_add3b_xor3b_wx117 = multm_reduce_mulb0_sq118 ^ multm_reduce_mulb0_cq117;
  assign multm_reduce_mulb0_add3b_xor3b_wx118 = multm_reduce_mulb0_sq119 ^ multm_reduce_mulb0_cq118;
  assign multm_reduce_mulb0_add3b_xor3b_wx120 = multm_reduce_mulb0_sq121 ^ multm_reduce_mulb0_cq120;
  assign multm_reduce_mulb0_add3b_xor3b_wx122 = multm_reduce_mulb0_sq123 ^ multm_reduce_mulb0_cq122;
  assign multm_reduce_mulb0_add3b_xor3b_wx123 = multm_reduce_mulb0_sq124 ^ multm_reduce_mulb0_cq123;
  assign multm_reduce_mulb0_add3b_xor3b_wx127 = multm_reduce_mulb0_sq128 ^ multm_reduce_mulb0_cq127;
  assign multm_reduce_mulb0_add3b_xor3b_wx128 = multm_reduce_mulb0_sq129 ^ multm_reduce_mulb0_cq128;
  assign multm_reduce_mulb0_add3b_xor3b_wx131 = multm_reduce_mulb0_sq132 ^ multm_reduce_mulb0_cq131;
  assign multm_reduce_mulb0_add3b_xor3b_wx134 = multm_reduce_mulb0_sq135 ^ multm_reduce_mulb0_cq134;
  assign multm_reduce_mulb0_add3b_xor3b_wx135 = multm_reduce_mulb0_sq136 ^ multm_reduce_mulb0_cq135;
  assign multm_reduce_mulb0_add3b_xor3b_wx136 = multm_reduce_mulb0_sq137 ^ multm_reduce_mulb0_cq136;
  assign multm_reduce_mulb0_add3b_xor3b_wx138 = multm_reduce_mulb0_sq139 ^ multm_reduce_mulb0_cq138;
  assign multm_reduce_mulb0_add3b_xor3b_wx140 = multm_reduce_mulb0_sq141 ^ multm_reduce_mulb0_cq140;
  assign multm_reduce_mulb0_add3b_xor3b_wx146 = multm_reduce_mulb0_sq147 ^ multm_reduce_mulb0_cq146;
  assign multm_reduce_mulb0_add3b_xor3b_wx147 = multm_reduce_mulb0_sq148 ^ multm_reduce_mulb0_cq147;
  assign multm_reduce_mulb0_add3b_xor3b_wx148 = multm_reduce_mulb0_sq149 ^ multm_reduce_mulb0_cq148;
  assign multm_reduce_mulb0_add3b_xor3b_wx149 = multm_reduce_mulb0_sq150 ^ multm_reduce_mulb0_cq149;
  assign multm_reduce_mulb0_add3b_xor3b_wx152 = multm_reduce_mulb0_sq153 ^ multm_reduce_mulb0_cq152;
  assign multm_reduce_mulb0_add3b_xor3b_wx153 = multm_reduce_mulb0_sq154 ^ multm_reduce_mulb0_cq153;
  assign multm_reduce_mulb0_add3b_xor3b_wx156 = multm_reduce_mulb0_sq157 ^ multm_reduce_mulb0_cq156;
  assign multm_reduce_mulb0_add3b_xor3b_wx157 = multm_reduce_mulb0_sq158 ^ multm_reduce_mulb0_cq157;
  assign multm_reduce_mulb0_add3b_xor3b_wx158 = multm_reduce_mulb0_sq159 ^ multm_reduce_mulb0_cq158;
  assign multm_reduce_mulb0_add3b_xor3b_wx159 = multm_reduce_mulb0_sq160 ^ multm_reduce_mulb0_cq159;
  assign multm_reduce_mulb0_add3b_xor3b_wx160 = multm_reduce_mulb0_sq161 ^ multm_reduce_mulb0_cq160;
  assign multm_reduce_mulb0_add3b_xor3b_wx162 = multm_reduce_mulb0_sq163 ^ multm_reduce_mulb0_cq162;
  assign multm_reduce_mulb0_add3b_xor3b_wx163 = multm_reduce_mulb0_sq164 ^ multm_reduce_mulb0_cq163;
  assign multm_reduce_mulb0_add3b_xor3b_wx168 = multm_reduce_mulb0_sq169 ^ multm_reduce_mulb0_cq168;
  assign multm_reduce_mulb0_add3b_xor3b_wx170 = multm_reduce_mulb0_sq171 ^ multm_reduce_mulb0_cq170;
  assign multm_reduce_mulb0_add3b_xor3b_wx171 = multm_reduce_mulb0_sq172 ^ multm_reduce_mulb0_cq171;
  assign multm_reduce_mulb0_add3b_xor3b_wx172 = multm_reduce_mulb0_sq173 ^ multm_reduce_mulb0_cq172;
  assign multm_reduce_mulb0_add3b_xor3b_wx173 = multm_reduce_mulb0_sq174 ^ multm_reduce_mulb0_cq173;
  assign multm_reduce_mulb0_add3b_xor3b_wx175 = multm_reduce_mulb0_sq176 ^ multm_reduce_mulb0_cq175;
  assign multm_reduce_mulb0_add3b_xor3b_wx177 = multm_reduce_mulb0_sq178 ^ multm_reduce_mulb0_cq177;
  assign multm_reduce_mulb0_add3b_xor3b_wx178 = multm_reduce_mulb0_sq179 ^ multm_reduce_mulb0_cq178;
  assign multm_reduce_mulb0_add3b_xor3b_wx181 = multm_reduce_mulb0_sq182 ^ multm_reduce_mulb0_cq181;
  assign multm_reduce_mulb0_add3b_xor3b_wx182 = multm_reduce_mulb0_sq183 ^ multm_reduce_mulb0_cq182;
  assign multm_reduce_mulb0_add3b_xor3b_wx183 = multm_reduce_mulb0_sq184 ^ multm_reduce_mulb0_cq183;
  assign multm_reduce_mulb0_cq0 = xn1 & multm_reduce_mulb0_cp0;
  assign multm_reduce_mulb0_cq1 = xn1 & multm_reduce_mulb0_cp1;
  assign multm_reduce_mulb0_cq2 = xn1 & multm_reduce_mulb0_cp2;
  assign multm_reduce_mulb0_cq3 = xn1 & multm_reduce_mulb0_cp3;
  assign multm_reduce_mulb0_cq4 = xn1 & multm_reduce_mulb0_cp4;
  assign multm_reduce_mulb0_cq5 = xn1 & multm_reduce_mulb0_cp5;
  assign multm_reduce_mulb0_cq6 = xn1 & multm_reduce_mulb0_cp6;
  assign multm_reduce_mulb0_cq7 = xn1 & multm_reduce_mulb0_cp7;
  assign multm_reduce_mulb0_cq8 = xn1 & multm_reduce_mulb0_cp8;
  assign multm_reduce_mulb0_cq9 = xn1 & multm_reduce_mulb0_cp9;
  assign multm_reduce_mulb0_cq10 = xn1 & multm_reduce_mulb0_cp10;
  assign multm_reduce_mulb0_cq11 = xn1 & multm_reduce_mulb0_cp11;
  assign multm_reduce_mulb0_cq12 = xn1 & multm_reduce_mulb0_cp12;
  assign multm_reduce_mulb0_cq13 = xn1 & multm_reduce_mulb0_cp13;
  assign multm_reduce_mulb0_cq14 = xn1 & multm_reduce_mulb0_cp14;
  assign multm_reduce_mulb0_cq15 = xn1 & multm_reduce_mulb0_cp15;
  assign multm_reduce_mulb0_cq16 = xn1 & multm_reduce_mulb0_cp16;
  assign multm_reduce_mulb0_cq17 = xn1 & multm_reduce_mulb0_cp17;
  assign multm_reduce_mulb0_cq18 = xn1 & multm_reduce_mulb0_cp18;
  assign multm_reduce_mulb0_cq19 = xn1 & multm_reduce_mulb0_cp19;
  assign multm_reduce_mulb0_cq20 = xn1 & multm_reduce_mulb0_cp20;
  assign multm_reduce_mulb0_cq21 = xn1 & multm_reduce_mulb0_cp21;
  assign multm_reduce_mulb0_cq22 = xn1 & multm_reduce_mulb0_cp22;
  assign multm_reduce_mulb0_cq23 = xn1 & multm_reduce_mulb0_cp23;
  assign multm_reduce_mulb0_cq24 = xn1 & multm_reduce_mulb0_cp24;
  assign multm_reduce_mulb0_cq25 = xn1 & multm_reduce_mulb0_cp25;
  assign multm_reduce_mulb0_cq26 = xn1 & multm_reduce_mulb0_cp26;
  assign multm_reduce_mulb0_cq27 = xn1 & multm_reduce_mulb0_cp27;
  assign multm_reduce_mulb0_cq28 = xn1 & multm_reduce_mulb0_cp28;
  assign multm_reduce_mulb0_cq29 = xn1 & multm_reduce_mulb0_cp29;
  assign multm_reduce_mulb0_cq30 = xn1 & multm_reduce_mulb0_cp30;
  assign multm_reduce_mulb0_cq31 = xn1 & multm_reduce_mulb0_cp31;
  assign multm_reduce_mulb0_cq32 = xn1 & multm_reduce_mulb0_cp32;
  assign multm_reduce_mulb0_cq33 = xn1 & multm_reduce_mulb0_cp33;
  assign multm_reduce_mulb0_cq34 = xn1 & multm_reduce_mulb0_cp34;
  assign multm_reduce_mulb0_cq35 = xn1 & multm_reduce_mulb0_cp35;
  assign multm_reduce_mulb0_cq36 = xn1 & multm_reduce_mulb0_cp36;
  assign multm_reduce_mulb0_cq37 = xn1 & multm_reduce_mulb0_cp37;
  assign multm_reduce_mulb0_cq38 = xn1 & multm_reduce_mulb0_cp38;
  assign multm_reduce_mulb0_cq39 = xn1 & multm_reduce_mulb0_cp39;
  assign multm_reduce_mulb0_cq40 = xn1 & multm_reduce_mulb0_cp40;
  assign multm_reduce_mulb0_cq41 = xn1 & multm_reduce_mulb0_cp41;
  assign multm_reduce_mulb0_cq42 = xn1 & multm_reduce_mulb0_cp42;
  assign multm_reduce_mulb0_cq43 = xn1 & multm_reduce_mulb0_cp43;
  assign multm_reduce_mulb0_cq44 = xn1 & multm_reduce_mulb0_cp44;
  assign multm_reduce_mulb0_cq45 = xn1 & multm_reduce_mulb0_cp45;
  assign multm_reduce_mulb0_cq46 = xn1 & multm_reduce_mulb0_cp46;
  assign multm_reduce_mulb0_cq47 = xn1 & multm_reduce_mulb0_cp47;
  assign multm_reduce_mulb0_cq48 = xn1 & multm_reduce_mulb0_cp48;
  assign multm_reduce_mulb0_cq49 = xn1 & multm_reduce_mulb0_cp49;
  assign multm_reduce_mulb0_cq50 = xn1 & multm_reduce_mulb0_cp50;
  assign multm_reduce_mulb0_cq51 = xn1 & multm_reduce_mulb0_cp51;
  assign multm_reduce_mulb0_cq52 = xn1 & multm_reduce_mulb0_cp52;
  assign multm_reduce_mulb0_cq53 = xn1 & multm_reduce_mulb0_cp53;
  assign multm_reduce_mulb0_cq54 = xn1 & multm_reduce_mulb0_cp54;
  assign multm_reduce_mulb0_cq55 = xn1 & multm_reduce_mulb0_cp55;
  assign multm_reduce_mulb0_cq56 = xn1 & multm_reduce_mulb0_cp56;
  assign multm_reduce_mulb0_cq57 = xn1 & multm_reduce_mulb0_cp57;
  assign multm_reduce_mulb0_cq58 = xn1 & multm_reduce_mulb0_cp58;
  assign multm_reduce_mulb0_cq59 = xn1 & multm_reduce_mulb0_cp59;
  assign multm_reduce_mulb0_cq60 = xn1 & multm_reduce_mulb0_cp60;
  assign multm_reduce_mulb0_cq61 = xn1 & multm_reduce_mulb0_cp61;
  assign multm_reduce_mulb0_cq62 = xn1 & multm_reduce_mulb0_cp62;
  assign multm_reduce_mulb0_cq63 = xn1 & multm_reduce_mulb0_cp63;
  assign multm_reduce_mulb0_cq64 = xn1 & multm_reduce_mulb0_cp64;
  assign multm_reduce_mulb0_cq65 = xn1 & multm_reduce_mulb0_cp65;
  assign multm_reduce_mulb0_cq66 = xn1 & multm_reduce_mulb0_cp66;
  assign multm_reduce_mulb0_cq67 = xn1 & multm_reduce_mulb0_cp67;
  assign multm_reduce_mulb0_cq68 = xn1 & multm_reduce_mulb0_cp68;
  assign multm_reduce_mulb0_cq69 = xn1 & multm_reduce_mulb0_cp69;
  assign multm_reduce_mulb0_cq70 = xn1 & multm_reduce_mulb0_cp70;
  assign multm_reduce_mulb0_cq71 = xn1 & multm_reduce_mulb0_cp71;
  assign multm_reduce_mulb0_cq72 = xn1 & multm_reduce_mulb0_cp72;
  assign multm_reduce_mulb0_cq73 = xn1 & multm_reduce_mulb0_cp73;
  assign multm_reduce_mulb0_cq74 = xn1 & multm_reduce_mulb0_cp74;
  assign multm_reduce_mulb0_cq75 = xn1 & multm_reduce_mulb0_cp75;
  assign multm_reduce_mulb0_cq76 = xn1 & multm_reduce_mulb0_cp76;
  assign multm_reduce_mulb0_cq77 = xn1 & multm_reduce_mulb0_cp77;
  assign multm_reduce_mulb0_cq78 = xn1 & multm_reduce_mulb0_cp78;
  assign multm_reduce_mulb0_cq79 = xn1 & multm_reduce_mulb0_cp79;
  assign multm_reduce_mulb0_cq80 = xn1 & multm_reduce_mulb0_cp80;
  assign multm_reduce_mulb0_cq81 = xn1 & multm_reduce_mulb0_cp81;
  assign multm_reduce_mulb0_cq82 = xn1 & multm_reduce_mulb0_cp82;
  assign multm_reduce_mulb0_cq83 = xn1 & multm_reduce_mulb0_cp83;
  assign multm_reduce_mulb0_cq84 = xn1 & multm_reduce_mulb0_cp84;
  assign multm_reduce_mulb0_cq85 = xn1 & multm_reduce_mulb0_cp85;
  assign multm_reduce_mulb0_cq86 = xn1 & multm_reduce_mulb0_cp86;
  assign multm_reduce_mulb0_cq87 = xn1 & multm_reduce_mulb0_cp87;
  assign multm_reduce_mulb0_cq88 = xn1 & multm_reduce_mulb0_cp88;
  assign multm_reduce_mulb0_cq89 = xn1 & multm_reduce_mulb0_cp89;
  assign multm_reduce_mulb0_cq90 = xn1 & multm_reduce_mulb0_cp90;
  assign multm_reduce_mulb0_cq91 = xn1 & multm_reduce_mulb0_cp91;
  assign multm_reduce_mulb0_cq92 = xn1 & multm_reduce_mulb0_cp92;
  assign multm_reduce_mulb0_cq93 = xn1 & multm_reduce_mulb0_cp93;
  assign multm_reduce_mulb0_cq94 = xn1 & multm_reduce_mulb0_cp94;
  assign multm_reduce_mulb0_cq95 = xn1 & multm_reduce_mulb0_cp95;
  assign multm_reduce_mulb0_cq96 = xn1 & multm_reduce_mulb0_cp96;
  assign multm_reduce_mulb0_cq97 = xn1 & multm_reduce_mulb0_cp97;
  assign multm_reduce_mulb0_cq98 = xn1 & multm_reduce_mulb0_cp98;
  assign multm_reduce_mulb0_cq99 = xn1 & multm_reduce_mulb0_cp99;
  assign multm_reduce_mulb0_cq100 = xn1 & multm_reduce_mulb0_cp100;
  assign multm_reduce_mulb0_cq101 = xn1 & multm_reduce_mulb0_cp101;
  assign multm_reduce_mulb0_cq102 = xn1 & multm_reduce_mulb0_cp102;
  assign multm_reduce_mulb0_cq103 = xn1 & multm_reduce_mulb0_cp103;
  assign multm_reduce_mulb0_cq104 = xn1 & multm_reduce_mulb0_cp104;
  assign multm_reduce_mulb0_cq105 = xn1 & multm_reduce_mulb0_cp105;
  assign multm_reduce_mulb0_cq106 = xn1 & multm_reduce_mulb0_cp106;
  assign multm_reduce_mulb0_cq107 = xn1 & multm_reduce_mulb0_cp107;
  assign multm_reduce_mulb0_cq108 = xn1 & multm_reduce_mulb0_cp108;
  assign multm_reduce_mulb0_cq109 = xn1 & multm_reduce_mulb0_cp109;
  assign multm_reduce_mulb0_cq110 = xn1 & multm_reduce_mulb0_cp110;
  assign multm_reduce_mulb0_cq111 = xn1 & multm_reduce_mulb0_cp111;
  assign multm_reduce_mulb0_cq112 = xn1 & multm_reduce_mulb0_cp112;
  assign multm_reduce_mulb0_cq113 = xn1 & multm_reduce_mulb0_cp113;
  assign multm_reduce_mulb0_cq114 = xn1 & multm_reduce_mulb0_cp114;
  assign multm_reduce_mulb0_cq115 = xn1 & multm_reduce_mulb0_cp115;
  assign multm_reduce_mulb0_cq116 = xn1 & multm_reduce_mulb0_cp116;
  assign multm_reduce_mulb0_cq117 = xn1 & multm_reduce_mulb0_cp117;
  assign multm_reduce_mulb0_cq118 = xn1 & multm_reduce_mulb0_cp118;
  assign multm_reduce_mulb0_cq119 = xn1 & multm_reduce_mulb0_cp119;
  assign multm_reduce_mulb0_cq120 = xn1 & multm_reduce_mulb0_cp120;
  assign multm_reduce_mulb0_cq121 = xn1 & multm_reduce_mulb0_cp121;
  assign multm_reduce_mulb0_cq122 = xn1 & multm_reduce_mulb0_cp122;
  assign multm_reduce_mulb0_cq123 = xn1 & multm_reduce_mulb0_cp123;
  assign multm_reduce_mulb0_cq124 = xn1 & multm_reduce_mulb0_cp124;
  assign multm_reduce_mulb0_cq125 = xn1 & multm_reduce_mulb0_cp125;
  assign multm_reduce_mulb0_cq126 = xn1 & multm_reduce_mulb0_cp126;
  assign multm_reduce_mulb0_cq127 = xn1 & multm_reduce_mulb0_cp127;
  assign multm_reduce_mulb0_cq128 = xn1 & multm_reduce_mulb0_cp128;
  assign multm_reduce_mulb0_cq129 = xn1 & multm_reduce_mulb0_cp129;
  assign multm_reduce_mulb0_cq130 = xn1 & multm_reduce_mulb0_cp130;
  assign multm_reduce_mulb0_cq131 = xn1 & multm_reduce_mulb0_cp131;
  assign multm_reduce_mulb0_cq132 = xn1 & multm_reduce_mulb0_cp132;
  assign multm_reduce_mulb0_cq133 = xn1 & multm_reduce_mulb0_cp133;
  assign multm_reduce_mulb0_cq134 = xn1 & multm_reduce_mulb0_cp134;
  assign multm_reduce_mulb0_cq135 = xn1 & multm_reduce_mulb0_cp135;
  assign multm_reduce_mulb0_cq136 = xn1 & multm_reduce_mulb0_cp136;
  assign multm_reduce_mulb0_cq137 = xn1 & multm_reduce_mulb0_cp137;
  assign multm_reduce_mulb0_cq138 = xn1 & multm_reduce_mulb0_cp138;
  assign multm_reduce_mulb0_cq139 = xn1 & multm_reduce_mulb0_cp139;
  assign multm_reduce_mulb0_cq140 = xn1 & multm_reduce_mulb0_cp140;
  assign multm_reduce_mulb0_cq141 = xn1 & multm_reduce_mulb0_cp141;
  assign multm_reduce_mulb0_cq142 = xn1 & multm_reduce_mulb0_cp142;
  assign multm_reduce_mulb0_cq143 = xn1 & multm_reduce_mulb0_cp143;
  assign multm_reduce_mulb0_cq144 = xn1 & multm_reduce_mulb0_cp144;
  assign multm_reduce_mulb0_cq145 = xn1 & multm_reduce_mulb0_cp145;
  assign multm_reduce_mulb0_cq146 = xn1 & multm_reduce_mulb0_cp146;
  assign multm_reduce_mulb0_cq147 = xn1 & multm_reduce_mulb0_cp147;
  assign multm_reduce_mulb0_cq148 = xn1 & multm_reduce_mulb0_cp148;
  assign multm_reduce_mulb0_cq149 = xn1 & multm_reduce_mulb0_cp149;
  assign multm_reduce_mulb0_cq150 = xn1 & multm_reduce_mulb0_cp150;
  assign multm_reduce_mulb0_cq151 = xn1 & multm_reduce_mulb0_cp151;
  assign multm_reduce_mulb0_cq152 = xn1 & multm_reduce_mulb0_cp152;
  assign multm_reduce_mulb0_cq153 = xn1 & multm_reduce_mulb0_cp153;
  assign multm_reduce_mulb0_cq154 = xn1 & multm_reduce_mulb0_cp154;
  assign multm_reduce_mulb0_cq155 = xn1 & multm_reduce_mulb0_cp155;
  assign multm_reduce_mulb0_cq156 = xn1 & multm_reduce_mulb0_cp156;
  assign multm_reduce_mulb0_cq157 = xn1 & multm_reduce_mulb0_cp157;
  assign multm_reduce_mulb0_cq158 = xn1 & multm_reduce_mulb0_cp158;
  assign multm_reduce_mulb0_cq159 = xn1 & multm_reduce_mulb0_cp159;
  assign multm_reduce_mulb0_cq160 = xn1 & multm_reduce_mulb0_cp160;
  assign multm_reduce_mulb0_cq161 = xn1 & multm_reduce_mulb0_cp161;
  assign multm_reduce_mulb0_cq162 = xn1 & multm_reduce_mulb0_cp162;
  assign multm_reduce_mulb0_cq163 = xn1 & multm_reduce_mulb0_cp163;
  assign multm_reduce_mulb0_cq164 = xn1 & multm_reduce_mulb0_cp164;
  assign multm_reduce_mulb0_cq165 = xn1 & multm_reduce_mulb0_cp165;
  assign multm_reduce_mulb0_cq166 = xn1 & multm_reduce_mulb0_cp166;
  assign multm_reduce_mulb0_cq167 = xn1 & multm_reduce_mulb0_cp167;
  assign multm_reduce_mulb0_cq168 = xn1 & multm_reduce_mulb0_cp168;
  assign multm_reduce_mulb0_cq169 = xn1 & multm_reduce_mulb0_cp169;
  assign multm_reduce_mulb0_cq170 = xn1 & multm_reduce_mulb0_cp170;
  assign multm_reduce_mulb0_cq171 = xn1 & multm_reduce_mulb0_cp171;
  assign multm_reduce_mulb0_cq172 = xn1 & multm_reduce_mulb0_cp172;
  assign multm_reduce_mulb0_cq173 = xn1 & multm_reduce_mulb0_cp173;
  assign multm_reduce_mulb0_cq174 = xn1 & multm_reduce_mulb0_cp174;
  assign multm_reduce_mulb0_cq175 = xn1 & multm_reduce_mulb0_cp175;
  assign multm_reduce_mulb0_cq176 = xn1 & multm_reduce_mulb0_cp176;
  assign multm_reduce_mulb0_cq177 = xn1 & multm_reduce_mulb0_cp177;
  assign multm_reduce_mulb0_cq178 = xn1 & multm_reduce_mulb0_cp178;
  assign multm_reduce_mulb0_cq179 = xn1 & multm_reduce_mulb0_cp179;
  assign multm_reduce_mulb0_cq180 = xn1 & multm_reduce_mulb0_cp180;
  assign multm_reduce_mulb0_cq181 = xn1 & multm_reduce_mulb0_cp181;
  assign multm_reduce_mulb0_cq182 = xn1 & multm_reduce_mulb0_cp182;
  assign multm_reduce_mulb0_cq183 = xn1 & multm_reduce_mulb0_cp183;
  assign multm_reduce_mulb0_cq184 = xn1 & multm_reduce_mulb0_cp184;
  assign multm_reduce_mulb0_pc0 = multm_reduce_mulb0_sq0 & multm_reduce_sa5;
  assign multm_reduce_mulb0_pc1 = multm_reduce_mulb0_sq1 & multm_reduce_mulb0_cq0;
  assign multm_reduce_mulb0_pc2 = multm_reduce_mulb0_sq2 & multm_reduce_mulb0_cq1;
  assign multm_reduce_mulb0_pc3 = multm_reduce_mulb0_add3b_maj3b_or3b_wx2 | multm_reduce_mulb0_add3b_maj3b_xy2;
  assign multm_reduce_mulb0_pc4 = multm_reduce_mulb0_sq4 & multm_reduce_mulb0_cq3;
  assign multm_reduce_mulb0_pc5 = multm_reduce_mulb0_add3b_maj3b_or3b_wx4 | multm_reduce_mulb0_add3b_maj3b_xy4;
  assign multm_reduce_mulb0_pc6 = multm_reduce_mulb0_sq6 & multm_reduce_mulb0_cq5;
  assign multm_reduce_mulb0_pc7 = multm_reduce_mulb0_sq7 & multm_reduce_mulb0_cq6;
  assign multm_reduce_mulb0_pc8 = multm_reduce_mulb0_sq8 & multm_reduce_mulb0_cq7;
  assign multm_reduce_mulb0_pc9 = multm_reduce_mulb0_add3b_maj3b_or3b_wx8 | multm_reduce_mulb0_add3b_maj3b_xy8;
  assign multm_reduce_mulb0_pc10 = multm_reduce_mulb0_add3b_maj3b_or3b_wx9 | multm_reduce_mulb0_add3b_maj3b_xy9;
  assign multm_reduce_mulb0_pc11 = multm_reduce_mulb0_sq11 & multm_reduce_mulb0_cq10;
  assign multm_reduce_mulb0_pc12 = multm_reduce_mulb0_sq12 & multm_reduce_mulb0_cq11;
  assign multm_reduce_mulb0_pc13 = multm_reduce_mulb0_add3b_maj3b_or3b_wx12 | multm_reduce_mulb0_add3b_maj3b_xy12;
  assign multm_reduce_mulb0_pc14 = multm_reduce_mulb0_sq14 & multm_reduce_mulb0_cq13;
  assign multm_reduce_mulb0_pc15 = multm_reduce_mulb0_sq15 & multm_reduce_mulb0_cq14;
  assign multm_reduce_mulb0_pc16 = multm_reduce_mulb0_add3b_maj3b_or3b_wx15 | multm_reduce_mulb0_add3b_maj3b_xy15;
  assign multm_reduce_mulb0_pc17 = multm_reduce_mulb0_add3b_maj3b_or3b_wx16 | multm_reduce_mulb0_add3b_maj3b_xy16;
  assign multm_reduce_mulb0_pc18 = multm_reduce_mulb0_add3b_maj3b_or3b_wx17 | multm_reduce_mulb0_add3b_maj3b_xy17;
  assign multm_reduce_mulb0_pc19 = multm_reduce_mulb0_add3b_maj3b_or3b_wx18 | multm_reduce_mulb0_add3b_maj3b_xy18;
  assign multm_reduce_mulb0_pc20 = multm_reduce_mulb0_add3b_maj3b_or3b_wx19 | multm_reduce_mulb0_add3b_maj3b_xy19;
  assign multm_reduce_mulb0_pc21 = multm_reduce_mulb0_add3b_maj3b_or3b_wx20 | multm_reduce_mulb0_add3b_maj3b_xy20;
  assign multm_reduce_mulb0_pc22 = multm_reduce_mulb0_sq22 & multm_reduce_mulb0_cq21;
  assign multm_reduce_mulb0_pc23 = multm_reduce_mulb0_sq23 & multm_reduce_mulb0_cq22;
  assign multm_reduce_mulb0_pc24 = multm_reduce_mulb0_sq24 & multm_reduce_mulb0_cq23;
  assign multm_reduce_mulb0_pc25 = multm_reduce_mulb0_sq25 & multm_reduce_mulb0_cq24;
  assign multm_reduce_mulb0_pc26 = multm_reduce_mulb0_add3b_maj3b_or3b_wx25 | multm_reduce_mulb0_add3b_maj3b_xy25;
  assign multm_reduce_mulb0_pc27 = multm_reduce_mulb0_add3b_maj3b_or3b_wx26 | multm_reduce_mulb0_add3b_maj3b_xy26;
  assign multm_reduce_mulb0_pc28 = multm_reduce_mulb0_add3b_maj3b_or3b_wx27 | multm_reduce_mulb0_add3b_maj3b_xy27;
  assign multm_reduce_mulb0_pc29 = multm_reduce_mulb0_sq29 & multm_reduce_mulb0_cq28;
  assign multm_reduce_mulb0_pc30 = multm_reduce_mulb0_add3b_maj3b_or3b_wx29 | multm_reduce_mulb0_add3b_maj3b_xy29;
  assign multm_reduce_mulb0_pc31 = multm_reduce_mulb0_add3b_maj3b_or3b_wx30 | multm_reduce_mulb0_add3b_maj3b_xy30;
  assign multm_reduce_mulb0_pc32 = multm_reduce_mulb0_sq32 & multm_reduce_mulb0_cq31;
  assign multm_reduce_mulb0_pc33 = multm_reduce_mulb0_sq33 & multm_reduce_mulb0_cq32;
  assign multm_reduce_mulb0_pc34 = multm_reduce_mulb0_add3b_maj3b_or3b_wx33 | multm_reduce_mulb0_add3b_maj3b_xy33;
  assign multm_reduce_mulb0_pc35 = multm_reduce_mulb0_sq35 & multm_reduce_mulb0_cq34;
  assign multm_reduce_mulb0_pc36 = multm_reduce_mulb0_sq36 & multm_reduce_mulb0_cq35;
  assign multm_reduce_mulb0_pc37 = multm_reduce_mulb0_sq37 & multm_reduce_mulb0_cq36;
  assign multm_reduce_mulb0_pc38 = multm_reduce_mulb0_add3b_maj3b_or3b_wx37 | multm_reduce_mulb0_add3b_maj3b_xy37;
  assign multm_reduce_mulb0_pc39 = multm_reduce_mulb0_sq39 & multm_reduce_mulb0_cq38;
  assign multm_reduce_mulb0_pc40 = multm_reduce_mulb0_sq40 & multm_reduce_mulb0_cq39;
  assign multm_reduce_mulb0_pc41 = multm_reduce_mulb0_add3b_maj3b_or3b_wx40 | multm_reduce_mulb0_add3b_maj3b_xy40;
  assign multm_reduce_mulb0_pc42 = multm_reduce_mulb0_sq42 & multm_reduce_mulb0_cq41;
  assign multm_reduce_mulb0_pc43 = multm_reduce_mulb0_add3b_maj3b_or3b_wx42 | multm_reduce_mulb0_add3b_maj3b_xy42;
  assign multm_reduce_mulb0_pc44 = multm_reduce_mulb0_sq44 & multm_reduce_mulb0_cq43;
  assign multm_reduce_mulb0_pc45 = multm_reduce_mulb0_add3b_maj3b_or3b_wx44 | multm_reduce_mulb0_add3b_maj3b_xy44;
  assign multm_reduce_mulb0_pc46 = multm_reduce_mulb0_add3b_maj3b_or3b_wx45 | multm_reduce_mulb0_add3b_maj3b_xy45;
  assign multm_reduce_mulb0_pc47 = multm_reduce_mulb0_add3b_maj3b_or3b_wx46 | multm_reduce_mulb0_add3b_maj3b_xy46;
  assign multm_reduce_mulb0_pc48 = multm_reduce_mulb0_sq48 & multm_reduce_mulb0_cq47;
  assign multm_reduce_mulb0_pc49 = multm_reduce_mulb0_add3b_maj3b_or3b_wx48 | multm_reduce_mulb0_add3b_maj3b_xy48;
  assign multm_reduce_mulb0_pc50 = multm_reduce_mulb0_sq50 & multm_reduce_mulb0_cq49;
  assign multm_reduce_mulb0_pc51 = multm_reduce_mulb0_add3b_maj3b_or3b_wx50 | multm_reduce_mulb0_add3b_maj3b_xy50;
  assign multm_reduce_mulb0_pc52 = multm_reduce_mulb0_add3b_maj3b_or3b_wx51 | multm_reduce_mulb0_add3b_maj3b_xy51;
  assign multm_reduce_mulb0_pc53 = multm_reduce_mulb0_add3b_maj3b_or3b_wx52 | multm_reduce_mulb0_add3b_maj3b_xy52;
  assign multm_reduce_mulb0_pc54 = multm_reduce_mulb0_add3b_maj3b_or3b_wx53 | multm_reduce_mulb0_add3b_maj3b_xy53;
  assign multm_reduce_mulb0_pc55 = multm_reduce_mulb0_add3b_maj3b_or3b_wx54 | multm_reduce_mulb0_add3b_maj3b_xy54;
  assign multm_reduce_mulb0_pc56 = multm_reduce_mulb0_sq56 & multm_reduce_mulb0_cq55;
  assign multm_reduce_mulb0_pc57 = multm_reduce_mulb0_add3b_maj3b_or3b_wx56 | multm_reduce_mulb0_add3b_maj3b_xy56;
  assign multm_reduce_mulb0_pc58 = multm_reduce_mulb0_add3b_maj3b_or3b_wx57 | multm_reduce_mulb0_add3b_maj3b_xy57;
  assign multm_reduce_mulb0_pc59 = multm_reduce_mulb0_add3b_maj3b_or3b_wx58 | multm_reduce_mulb0_add3b_maj3b_xy58;
  assign multm_reduce_mulb0_pc60 = multm_reduce_mulb0_sq60 & multm_reduce_mulb0_cq59;
  assign multm_reduce_mulb0_pc61 = multm_reduce_mulb0_add3b_maj3b_or3b_wx60 | multm_reduce_mulb0_add3b_maj3b_xy60;
  assign multm_reduce_mulb0_pc62 = multm_reduce_mulb0_add3b_maj3b_or3b_wx61 | multm_reduce_mulb0_add3b_maj3b_xy61;
  assign multm_reduce_mulb0_pc63 = multm_reduce_mulb0_add3b_maj3b_or3b_wx62 | multm_reduce_mulb0_add3b_maj3b_xy62;
  assign multm_reduce_mulb0_pc64 = multm_reduce_mulb0_add3b_maj3b_or3b_wx63 | multm_reduce_mulb0_add3b_maj3b_xy63;
  assign multm_reduce_mulb0_pc65 = multm_reduce_mulb0_sq65 & multm_reduce_mulb0_cq64;
  assign multm_reduce_mulb0_pc66 = multm_reduce_mulb0_add3b_maj3b_or3b_wx65 | multm_reduce_mulb0_add3b_maj3b_xy65;
  assign multm_reduce_mulb0_pc67 = multm_reduce_mulb0_add3b_maj3b_or3b_wx66 | multm_reduce_mulb0_add3b_maj3b_xy66;
  assign multm_reduce_mulb0_pc68 = multm_reduce_mulb0_add3b_maj3b_or3b_wx67 | multm_reduce_mulb0_add3b_maj3b_xy67;
  assign multm_reduce_mulb0_pc69 = multm_reduce_mulb0_sq69 & multm_reduce_mulb0_cq68;
  assign multm_reduce_mulb0_pc70 = multm_reduce_mulb0_add3b_maj3b_or3b_wx69 | multm_reduce_mulb0_add3b_maj3b_xy69;
  assign multm_reduce_mulb0_pc71 = multm_reduce_mulb0_sq71 & multm_reduce_mulb0_cq70;
  assign multm_reduce_mulb0_pc72 = multm_reduce_mulb0_sq72 & multm_reduce_mulb0_cq71;
  assign multm_reduce_mulb0_pc73 = multm_reduce_mulb0_add3b_maj3b_or3b_wx72 | multm_reduce_mulb0_add3b_maj3b_xy72;
  assign multm_reduce_mulb0_pc74 = multm_reduce_mulb0_add3b_maj3b_or3b_wx73 | multm_reduce_mulb0_add3b_maj3b_xy73;
  assign multm_reduce_mulb0_pc75 = multm_reduce_mulb0_sq75 & multm_reduce_mulb0_cq74;
  assign multm_reduce_mulb0_pc76 = multm_reduce_mulb0_sq76 & multm_reduce_mulb0_cq75;
  assign multm_reduce_mulb0_pc77 = multm_reduce_mulb0_add3b_maj3b_or3b_wx76 | multm_reduce_mulb0_add3b_maj3b_xy76;
  assign multm_reduce_mulb0_pc78 = multm_reduce_mulb0_sq78 & multm_reduce_mulb0_cq77;
  assign multm_reduce_mulb0_pc79 = multm_reduce_mulb0_add3b_maj3b_or3b_wx78 | multm_reduce_mulb0_add3b_maj3b_xy78;
  assign multm_reduce_mulb0_pc80 = multm_reduce_mulb0_sq80 & multm_reduce_mulb0_cq79;
  assign multm_reduce_mulb0_pc81 = multm_reduce_mulb0_add3b_maj3b_or3b_wx80 | multm_reduce_mulb0_add3b_maj3b_xy80;
  assign multm_reduce_mulb0_pc82 = multm_reduce_mulb0_sq82 & multm_reduce_mulb0_cq81;
  assign multm_reduce_mulb0_pc83 = multm_reduce_mulb0_add3b_maj3b_or3b_wx82 | multm_reduce_mulb0_add3b_maj3b_xy82;
  assign multm_reduce_mulb0_pc84 = multm_reduce_mulb0_add3b_maj3b_or3b_wx83 | multm_reduce_mulb0_add3b_maj3b_xy83;
  assign multm_reduce_mulb0_pc85 = multm_reduce_mulb0_add3b_maj3b_or3b_wx84 | multm_reduce_mulb0_add3b_maj3b_xy84;
  assign multm_reduce_mulb0_pc86 = multm_reduce_mulb0_sq86 & multm_reduce_mulb0_cq85;
  assign multm_reduce_mulb0_pc87 = multm_reduce_mulb0_sq87 & multm_reduce_mulb0_cq86;
  assign multm_reduce_mulb0_pc88 = multm_reduce_mulb0_add3b_maj3b_or3b_wx87 | multm_reduce_mulb0_add3b_maj3b_xy87;
  assign multm_reduce_mulb0_pc89 = multm_reduce_mulb0_sq89 & multm_reduce_mulb0_cq88;
  assign multm_reduce_mulb0_pc90 = multm_reduce_mulb0_sq90 & multm_reduce_mulb0_cq89;
  assign multm_reduce_mulb0_pc91 = multm_reduce_mulb0_sq91 & multm_reduce_mulb0_cq90;
  assign multm_reduce_mulb0_pc92 = multm_reduce_mulb0_add3b_maj3b_or3b_wx91 | multm_reduce_mulb0_add3b_maj3b_xy91;
  assign multm_reduce_mulb0_pc93 = multm_reduce_mulb0_add3b_maj3b_or3b_wx92 | multm_reduce_mulb0_add3b_maj3b_xy92;
  assign multm_reduce_mulb0_pc94 = multm_reduce_mulb0_sq94 & multm_reduce_mulb0_cq93;
  assign multm_reduce_mulb0_pc95 = multm_reduce_mulb0_sq95 & multm_reduce_mulb0_cq94;
  assign multm_reduce_mulb0_pc96 = multm_reduce_mulb0_add3b_maj3b_or3b_wx95 | multm_reduce_mulb0_add3b_maj3b_xy95;
  assign multm_reduce_mulb0_pc97 = multm_reduce_mulb0_sq97 & multm_reduce_mulb0_cq96;
  assign multm_reduce_mulb0_pc98 = multm_reduce_mulb0_sq98 & multm_reduce_mulb0_cq97;
  assign multm_reduce_mulb0_pc99 = multm_reduce_mulb0_sq99 & multm_reduce_mulb0_cq98;
  assign multm_reduce_mulb0_pc100 = multm_reduce_mulb0_sq100 & multm_reduce_mulb0_cq99;
  assign multm_reduce_mulb0_pc101 = multm_reduce_mulb0_sq101 & multm_reduce_mulb0_cq100;
  assign multm_reduce_mulb0_pc102 = multm_reduce_mulb0_sq102 & multm_reduce_mulb0_cq101;
  assign multm_reduce_mulb0_pc103 = multm_reduce_mulb0_add3b_maj3b_or3b_wx102 | multm_reduce_mulb0_add3b_maj3b_xy102;
  assign multm_reduce_mulb0_pc104 = multm_reduce_mulb0_add3b_maj3b_or3b_wx103 | multm_reduce_mulb0_add3b_maj3b_xy103;
  assign multm_reduce_mulb0_pc105 = multm_reduce_mulb0_sq105 & multm_reduce_mulb0_cq104;
  assign multm_reduce_mulb0_pc106 = multm_reduce_mulb0_add3b_maj3b_or3b_wx105 | multm_reduce_mulb0_add3b_maj3b_xy105;
  assign multm_reduce_mulb0_pc107 = multm_reduce_mulb0_sq107 & multm_reduce_mulb0_cq106;
  assign multm_reduce_mulb0_pc108 = multm_reduce_mulb0_sq108 & multm_reduce_mulb0_cq107;
  assign multm_reduce_mulb0_pc109 = multm_reduce_mulb0_sq109 & multm_reduce_mulb0_cq108;
  assign multm_reduce_mulb0_pc110 = multm_reduce_mulb0_add3b_maj3b_or3b_wx109 | multm_reduce_mulb0_add3b_maj3b_xy109;
  assign multm_reduce_mulb0_pc111 = multm_reduce_mulb0_add3b_maj3b_or3b_wx110 | multm_reduce_mulb0_add3b_maj3b_xy110;
  assign multm_reduce_mulb0_pc112 = multm_reduce_mulb0_sq112 & multm_reduce_mulb0_cq111;
  assign multm_reduce_mulb0_pc113 = multm_reduce_mulb0_sq113 & multm_reduce_mulb0_cq112;
  assign multm_reduce_mulb0_pc114 = multm_reduce_mulb0_sq114 & multm_reduce_mulb0_cq113;
  assign multm_reduce_mulb0_pc115 = multm_reduce_mulb0_add3b_maj3b_or3b_wx114 | multm_reduce_mulb0_add3b_maj3b_xy114;
  assign multm_reduce_mulb0_pc116 = multm_reduce_mulb0_sq116 & multm_reduce_mulb0_cq115;
  assign multm_reduce_mulb0_pc117 = multm_reduce_mulb0_sq117 & multm_reduce_mulb0_cq116;
  assign multm_reduce_mulb0_pc118 = multm_reduce_mulb0_add3b_maj3b_or3b_wx117 | multm_reduce_mulb0_add3b_maj3b_xy117;
  assign multm_reduce_mulb0_pc119 = multm_reduce_mulb0_add3b_maj3b_or3b_wx118 | multm_reduce_mulb0_add3b_maj3b_xy118;
  assign multm_reduce_mulb0_pc120 = multm_reduce_mulb0_sq120 & multm_reduce_mulb0_cq119;
  assign multm_reduce_mulb0_pc121 = multm_reduce_mulb0_add3b_maj3b_or3b_wx120 | multm_reduce_mulb0_add3b_maj3b_xy120;
  assign multm_reduce_mulb0_pc122 = multm_reduce_mulb0_sq122 & multm_reduce_mulb0_cq121;
  assign multm_reduce_mulb0_pc123 = multm_reduce_mulb0_add3b_maj3b_or3b_wx122 | multm_reduce_mulb0_add3b_maj3b_xy122;
  assign multm_reduce_mulb0_pc124 = multm_reduce_mulb0_add3b_maj3b_or3b_wx123 | multm_reduce_mulb0_add3b_maj3b_xy123;
  assign multm_reduce_mulb0_pc125 = multm_reduce_mulb0_sq125 & multm_reduce_mulb0_cq124;
  assign multm_reduce_mulb0_pc126 = multm_reduce_mulb0_sq126 & multm_reduce_mulb0_cq125;
  assign multm_reduce_mulb0_pc127 = multm_reduce_mulb0_sq127 & multm_reduce_mulb0_cq126;
  assign multm_reduce_mulb0_pc128 = multm_reduce_mulb0_add3b_maj3b_or3b_wx127 | multm_reduce_mulb0_add3b_maj3b_xy127;
  assign multm_reduce_mulb0_pc129 = multm_reduce_mulb0_add3b_maj3b_or3b_wx128 | multm_reduce_mulb0_add3b_maj3b_xy128;
  assign multm_reduce_mulb0_pc130 = multm_reduce_mulb0_sq130 & multm_reduce_mulb0_cq129;
  assign multm_reduce_mulb0_pc131 = multm_reduce_mulb0_sq131 & multm_reduce_mulb0_cq130;
  assign multm_reduce_mulb0_pc132 = multm_reduce_mulb0_add3b_maj3b_or3b_wx131 | multm_reduce_mulb0_add3b_maj3b_xy131;
  assign multm_reduce_mulb0_pc133 = multm_reduce_mulb0_sq133 & multm_reduce_mulb0_cq132;
  assign multm_reduce_mulb0_pc134 = multm_reduce_mulb0_sq134 & multm_reduce_mulb0_cq133;
  assign multm_reduce_mulb0_pc135 = multm_reduce_mulb0_add3b_maj3b_or3b_wx134 | multm_reduce_mulb0_add3b_maj3b_xy134;
  assign multm_reduce_mulb0_pc136 = multm_reduce_mulb0_add3b_maj3b_or3b_wx135 | multm_reduce_mulb0_add3b_maj3b_xy135;
  assign multm_reduce_mulb0_pc137 = multm_reduce_mulb0_add3b_maj3b_or3b_wx136 | multm_reduce_mulb0_add3b_maj3b_xy136;
  assign multm_reduce_mulb0_pc138 = multm_reduce_mulb0_sq138 & multm_reduce_mulb0_cq137;
  assign multm_reduce_mulb0_pc139 = multm_reduce_mulb0_add3b_maj3b_or3b_wx138 | multm_reduce_mulb0_add3b_maj3b_xy138;
  assign multm_reduce_mulb0_pc140 = multm_reduce_mulb0_sq140 & multm_reduce_mulb0_cq139;
  assign multm_reduce_mulb0_pc141 = multm_reduce_mulb0_add3b_maj3b_or3b_wx140 | multm_reduce_mulb0_add3b_maj3b_xy140;
  assign multm_reduce_mulb0_pc142 = multm_reduce_mulb0_sq142 & multm_reduce_mulb0_cq141;
  assign multm_reduce_mulb0_pc143 = multm_reduce_mulb0_sq143 & multm_reduce_mulb0_cq142;
  assign multm_reduce_mulb0_pc144 = multm_reduce_mulb0_sq144 & multm_reduce_mulb0_cq143;
  assign multm_reduce_mulb0_pc145 = multm_reduce_mulb0_sq145 & multm_reduce_mulb0_cq144;
  assign multm_reduce_mulb0_pc146 = multm_reduce_mulb0_sq146 & multm_reduce_mulb0_cq145;
  assign multm_reduce_mulb0_pc147 = multm_reduce_mulb0_add3b_maj3b_or3b_wx146 | multm_reduce_mulb0_add3b_maj3b_xy146;
  assign multm_reduce_mulb0_pc148 = multm_reduce_mulb0_add3b_maj3b_or3b_wx147 | multm_reduce_mulb0_add3b_maj3b_xy147;
  assign multm_reduce_mulb0_pc149 = multm_reduce_mulb0_add3b_maj3b_or3b_wx148 | multm_reduce_mulb0_add3b_maj3b_xy148;
  assign multm_reduce_mulb0_pc150 = multm_reduce_mulb0_add3b_maj3b_or3b_wx149 | multm_reduce_mulb0_add3b_maj3b_xy149;
  assign multm_reduce_mulb0_pc151 = multm_reduce_mulb0_sq151 & multm_reduce_mulb0_cq150;
  assign multm_reduce_mulb0_pc152 = multm_reduce_mulb0_sq152 & multm_reduce_mulb0_cq151;
  assign multm_reduce_mulb0_pc153 = multm_reduce_mulb0_add3b_maj3b_or3b_wx152 | multm_reduce_mulb0_add3b_maj3b_xy152;
  assign multm_reduce_mulb0_pc154 = multm_reduce_mulb0_add3b_maj3b_or3b_wx153 | multm_reduce_mulb0_add3b_maj3b_xy153;
  assign multm_reduce_mulb0_pc155 = multm_reduce_mulb0_sq155 & multm_reduce_mulb0_cq154;
  assign multm_reduce_mulb0_pc156 = multm_reduce_mulb0_sq156 & multm_reduce_mulb0_cq155;
  assign multm_reduce_mulb0_pc157 = multm_reduce_mulb0_add3b_maj3b_or3b_wx156 | multm_reduce_mulb0_add3b_maj3b_xy156;
  assign multm_reduce_mulb0_pc158 = multm_reduce_mulb0_add3b_maj3b_or3b_wx157 | multm_reduce_mulb0_add3b_maj3b_xy157;
  assign multm_reduce_mulb0_pc159 = multm_reduce_mulb0_add3b_maj3b_or3b_wx158 | multm_reduce_mulb0_add3b_maj3b_xy158;
  assign multm_reduce_mulb0_pc160 = multm_reduce_mulb0_add3b_maj3b_or3b_wx159 | multm_reduce_mulb0_add3b_maj3b_xy159;
  assign multm_reduce_mulb0_pc161 = multm_reduce_mulb0_add3b_maj3b_or3b_wx160 | multm_reduce_mulb0_add3b_maj3b_xy160;
  assign multm_reduce_mulb0_pc162 = multm_reduce_mulb0_sq162 & multm_reduce_mulb0_cq161;
  assign multm_reduce_mulb0_pc163 = multm_reduce_mulb0_add3b_maj3b_or3b_wx162 | multm_reduce_mulb0_add3b_maj3b_xy162;
  assign multm_reduce_mulb0_pc164 = multm_reduce_mulb0_add3b_maj3b_or3b_wx163 | multm_reduce_mulb0_add3b_maj3b_xy163;
  assign multm_reduce_mulb0_pc165 = multm_reduce_mulb0_sq165 & multm_reduce_mulb0_cq164;
  assign multm_reduce_mulb0_pc166 = multm_reduce_mulb0_sq166 & multm_reduce_mulb0_cq165;
  assign multm_reduce_mulb0_pc167 = multm_reduce_mulb0_sq167 & multm_reduce_mulb0_cq166;
  assign multm_reduce_mulb0_pc168 = multm_reduce_mulb0_sq168 & multm_reduce_mulb0_cq167;
  assign multm_reduce_mulb0_pc169 = multm_reduce_mulb0_add3b_maj3b_or3b_wx168 | multm_reduce_mulb0_add3b_maj3b_xy168;
  assign multm_reduce_mulb0_pc170 = multm_reduce_mulb0_sq170 & multm_reduce_mulb0_cq169;
  assign multm_reduce_mulb0_pc171 = multm_reduce_mulb0_add3b_maj3b_or3b_wx170 | multm_reduce_mulb0_add3b_maj3b_xy170;
  assign multm_reduce_mulb0_pc172 = multm_reduce_mulb0_add3b_maj3b_or3b_wx171 | multm_reduce_mulb0_add3b_maj3b_xy171;
  assign multm_reduce_mulb0_pc173 = multm_reduce_mulb0_add3b_maj3b_or3b_wx172 | multm_reduce_mulb0_add3b_maj3b_xy172;
  assign multm_reduce_mulb0_pc174 = multm_reduce_mulb0_add3b_maj3b_or3b_wx173 | multm_reduce_mulb0_add3b_maj3b_xy173;
  assign multm_reduce_mulb0_pc175 = multm_reduce_mulb0_sq175 & multm_reduce_mulb0_cq174;
  assign multm_reduce_mulb0_pc176 = multm_reduce_mulb0_add3b_maj3b_or3b_wx175 | multm_reduce_mulb0_add3b_maj3b_xy175;
  assign multm_reduce_mulb0_pc177 = multm_reduce_mulb0_sq177 & multm_reduce_mulb0_cq176;
  assign multm_reduce_mulb0_pc178 = multm_reduce_mulb0_add3b_maj3b_or3b_wx177 | multm_reduce_mulb0_add3b_maj3b_xy177;
  assign multm_reduce_mulb0_pc179 = multm_reduce_mulb0_add3b_maj3b_or3b_wx178 | multm_reduce_mulb0_add3b_maj3b_xy178;
  assign multm_reduce_mulb0_pc180 = multm_reduce_mulb0_sq180 & multm_reduce_mulb0_cq179;
  assign multm_reduce_mulb0_pc181 = multm_reduce_mulb0_sq181 & multm_reduce_mulb0_cq180;
  assign multm_reduce_mulb0_pc182 = multm_reduce_mulb0_add3b_maj3b_or3b_wx181 | multm_reduce_mulb0_add3b_maj3b_xy181;
  assign multm_reduce_mulb0_pc183 = multm_reduce_mulb0_add3b_maj3b_or3b_wx182 | multm_reduce_mulb0_add3b_maj3b_xy182;
  assign multm_reduce_mulb0_pc184 = multm_reduce_mulb0_add3b_maj3b_or3b_wx183 | multm_reduce_mulb0_add3b_maj3b_xy183;
  assign multm_reduce_mulb0_ps0 = multm_reduce_mulb0_sq1 ^ multm_reduce_mulb0_cq0;
  assign multm_reduce_mulb0_ps1 = multm_reduce_mulb0_sq2 ^ multm_reduce_mulb0_cq1;
  assign multm_reduce_mulb0_ps2 = multm_reduce_mulb0_add3b_xor3b_wx2 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps3 = multm_reduce_mulb0_sq4 ^ multm_reduce_mulb0_cq3;
  assign multm_reduce_mulb0_ps4 = multm_reduce_mulb0_add3b_xor3b_wx4 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps5 = multm_reduce_mulb0_sq6 ^ multm_reduce_mulb0_cq5;
  assign multm_reduce_mulb0_ps6 = multm_reduce_mulb0_sq7 ^ multm_reduce_mulb0_cq6;
  assign multm_reduce_mulb0_ps7 = multm_reduce_mulb0_sq8 ^ multm_reduce_mulb0_cq7;
  assign multm_reduce_mulb0_ps8 = multm_reduce_mulb0_add3b_xor3b_wx8 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps9 = multm_reduce_mulb0_add3b_xor3b_wx9 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps10 = multm_reduce_mulb0_sq11 ^ multm_reduce_mulb0_cq10;
  assign multm_reduce_mulb0_ps11 = multm_reduce_mulb0_sq12 ^ multm_reduce_mulb0_cq11;
  assign multm_reduce_mulb0_ps12 = multm_reduce_mulb0_add3b_xor3b_wx12 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps13 = multm_reduce_mulb0_sq14 ^ multm_reduce_mulb0_cq13;
  assign multm_reduce_mulb0_ps14 = multm_reduce_mulb0_sq15 ^ multm_reduce_mulb0_cq14;
  assign multm_reduce_mulb0_ps15 = multm_reduce_mulb0_add3b_xor3b_wx15 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps16 = multm_reduce_mulb0_add3b_xor3b_wx16 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps17 = multm_reduce_mulb0_add3b_xor3b_wx17 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps18 = multm_reduce_mulb0_add3b_xor3b_wx18 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps19 = multm_reduce_mulb0_add3b_xor3b_wx19 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps20 = multm_reduce_mulb0_add3b_xor3b_wx20 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps21 = multm_reduce_mulb0_sq22 ^ multm_reduce_mulb0_cq21;
  assign multm_reduce_mulb0_ps22 = multm_reduce_mulb0_sq23 ^ multm_reduce_mulb0_cq22;
  assign multm_reduce_mulb0_ps23 = multm_reduce_mulb0_sq24 ^ multm_reduce_mulb0_cq23;
  assign multm_reduce_mulb0_ps24 = multm_reduce_mulb0_sq25 ^ multm_reduce_mulb0_cq24;
  assign multm_reduce_mulb0_ps25 = multm_reduce_mulb0_add3b_xor3b_wx25 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps26 = multm_reduce_mulb0_add3b_xor3b_wx26 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps27 = multm_reduce_mulb0_add3b_xor3b_wx27 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps28 = multm_reduce_mulb0_sq29 ^ multm_reduce_mulb0_cq28;
  assign multm_reduce_mulb0_ps29 = multm_reduce_mulb0_add3b_xor3b_wx29 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps30 = multm_reduce_mulb0_add3b_xor3b_wx30 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps31 = multm_reduce_mulb0_sq32 ^ multm_reduce_mulb0_cq31;
  assign multm_reduce_mulb0_ps32 = multm_reduce_mulb0_sq33 ^ multm_reduce_mulb0_cq32;
  assign multm_reduce_mulb0_ps33 = multm_reduce_mulb0_add3b_xor3b_wx33 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps34 = multm_reduce_mulb0_sq35 ^ multm_reduce_mulb0_cq34;
  assign multm_reduce_mulb0_ps35 = multm_reduce_mulb0_sq36 ^ multm_reduce_mulb0_cq35;
  assign multm_reduce_mulb0_ps36 = multm_reduce_mulb0_sq37 ^ multm_reduce_mulb0_cq36;
  assign multm_reduce_mulb0_ps37 = multm_reduce_mulb0_add3b_xor3b_wx37 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps38 = multm_reduce_mulb0_sq39 ^ multm_reduce_mulb0_cq38;
  assign multm_reduce_mulb0_ps39 = multm_reduce_mulb0_sq40 ^ multm_reduce_mulb0_cq39;
  assign multm_reduce_mulb0_ps40 = multm_reduce_mulb0_add3b_xor3b_wx40 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps41 = multm_reduce_mulb0_sq42 ^ multm_reduce_mulb0_cq41;
  assign multm_reduce_mulb0_ps42 = multm_reduce_mulb0_add3b_xor3b_wx42 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps43 = multm_reduce_mulb0_sq44 ^ multm_reduce_mulb0_cq43;
  assign multm_reduce_mulb0_ps44 = multm_reduce_mulb0_add3b_xor3b_wx44 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps45 = multm_reduce_mulb0_add3b_xor3b_wx45 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps46 = multm_reduce_mulb0_add3b_xor3b_wx46 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps47 = multm_reduce_mulb0_sq48 ^ multm_reduce_mulb0_cq47;
  assign multm_reduce_mulb0_ps48 = multm_reduce_mulb0_add3b_xor3b_wx48 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps49 = multm_reduce_mulb0_sq50 ^ multm_reduce_mulb0_cq49;
  assign multm_reduce_mulb0_ps50 = multm_reduce_mulb0_add3b_xor3b_wx50 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps51 = multm_reduce_mulb0_add3b_xor3b_wx51 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps52 = multm_reduce_mulb0_add3b_xor3b_wx52 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps53 = multm_reduce_mulb0_add3b_xor3b_wx53 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps54 = multm_reduce_mulb0_add3b_xor3b_wx54 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps55 = multm_reduce_mulb0_sq56 ^ multm_reduce_mulb0_cq55;
  assign multm_reduce_mulb0_ps56 = multm_reduce_mulb0_add3b_xor3b_wx56 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps57 = multm_reduce_mulb0_add3b_xor3b_wx57 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps58 = multm_reduce_mulb0_add3b_xor3b_wx58 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps59 = multm_reduce_mulb0_sq60 ^ multm_reduce_mulb0_cq59;
  assign multm_reduce_mulb0_ps60 = multm_reduce_mulb0_add3b_xor3b_wx60 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps61 = multm_reduce_mulb0_add3b_xor3b_wx61 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps62 = multm_reduce_mulb0_add3b_xor3b_wx62 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps63 = multm_reduce_mulb0_add3b_xor3b_wx63 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps64 = multm_reduce_mulb0_sq65 ^ multm_reduce_mulb0_cq64;
  assign multm_reduce_mulb0_ps65 = multm_reduce_mulb0_add3b_xor3b_wx65 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps66 = multm_reduce_mulb0_add3b_xor3b_wx66 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps67 = multm_reduce_mulb0_add3b_xor3b_wx67 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps68 = multm_reduce_mulb0_sq69 ^ multm_reduce_mulb0_cq68;
  assign multm_reduce_mulb0_ps69 = multm_reduce_mulb0_add3b_xor3b_wx69 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps70 = multm_reduce_mulb0_sq71 ^ multm_reduce_mulb0_cq70;
  assign multm_reduce_mulb0_ps71 = multm_reduce_mulb0_sq72 ^ multm_reduce_mulb0_cq71;
  assign multm_reduce_mulb0_ps72 = multm_reduce_mulb0_add3b_xor3b_wx72 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps73 = multm_reduce_mulb0_add3b_xor3b_wx73 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps74 = multm_reduce_mulb0_sq75 ^ multm_reduce_mulb0_cq74;
  assign multm_reduce_mulb0_ps75 = multm_reduce_mulb0_sq76 ^ multm_reduce_mulb0_cq75;
  assign multm_reduce_mulb0_ps76 = multm_reduce_mulb0_add3b_xor3b_wx76 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps77 = multm_reduce_mulb0_sq78 ^ multm_reduce_mulb0_cq77;
  assign multm_reduce_mulb0_ps78 = multm_reduce_mulb0_add3b_xor3b_wx78 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps79 = multm_reduce_mulb0_sq80 ^ multm_reduce_mulb0_cq79;
  assign multm_reduce_mulb0_ps80 = multm_reduce_mulb0_add3b_xor3b_wx80 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps81 = multm_reduce_mulb0_sq82 ^ multm_reduce_mulb0_cq81;
  assign multm_reduce_mulb0_ps82 = multm_reduce_mulb0_add3b_xor3b_wx82 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps83 = multm_reduce_mulb0_add3b_xor3b_wx83 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps84 = multm_reduce_mulb0_add3b_xor3b_wx84 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps85 = multm_reduce_mulb0_sq86 ^ multm_reduce_mulb0_cq85;
  assign multm_reduce_mulb0_ps86 = multm_reduce_mulb0_sq87 ^ multm_reduce_mulb0_cq86;
  assign multm_reduce_mulb0_ps87 = multm_reduce_mulb0_add3b_xor3b_wx87 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps88 = multm_reduce_mulb0_sq89 ^ multm_reduce_mulb0_cq88;
  assign multm_reduce_mulb0_ps89 = multm_reduce_mulb0_sq90 ^ multm_reduce_mulb0_cq89;
  assign multm_reduce_mulb0_ps90 = multm_reduce_mulb0_sq91 ^ multm_reduce_mulb0_cq90;
  assign multm_reduce_mulb0_ps91 = multm_reduce_mulb0_add3b_xor3b_wx91 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps92 = multm_reduce_mulb0_add3b_xor3b_wx92 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps93 = multm_reduce_mulb0_sq94 ^ multm_reduce_mulb0_cq93;
  assign multm_reduce_mulb0_ps94 = multm_reduce_mulb0_sq95 ^ multm_reduce_mulb0_cq94;
  assign multm_reduce_mulb0_ps95 = multm_reduce_mulb0_add3b_xor3b_wx95 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps96 = multm_reduce_mulb0_sq97 ^ multm_reduce_mulb0_cq96;
  assign multm_reduce_mulb0_ps97 = multm_reduce_mulb0_sq98 ^ multm_reduce_mulb0_cq97;
  assign multm_reduce_mulb0_ps98 = multm_reduce_mulb0_sq99 ^ multm_reduce_mulb0_cq98;
  assign multm_reduce_mulb0_ps99 = multm_reduce_mulb0_sq100 ^ multm_reduce_mulb0_cq99;
  assign multm_reduce_mulb0_ps100 = multm_reduce_mulb0_sq101 ^ multm_reduce_mulb0_cq100;
  assign multm_reduce_mulb0_ps101 = multm_reduce_mulb0_sq102 ^ multm_reduce_mulb0_cq101;
  assign multm_reduce_mulb0_ps102 = multm_reduce_mulb0_add3b_xor3b_wx102 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps103 = multm_reduce_mulb0_add3b_xor3b_wx103 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps104 = multm_reduce_mulb0_sq105 ^ multm_reduce_mulb0_cq104;
  assign multm_reduce_mulb0_ps105 = multm_reduce_mulb0_add3b_xor3b_wx105 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps106 = multm_reduce_mulb0_sq107 ^ multm_reduce_mulb0_cq106;
  assign multm_reduce_mulb0_ps107 = multm_reduce_mulb0_sq108 ^ multm_reduce_mulb0_cq107;
  assign multm_reduce_mulb0_ps108 = multm_reduce_mulb0_sq109 ^ multm_reduce_mulb0_cq108;
  assign multm_reduce_mulb0_ps109 = multm_reduce_mulb0_add3b_xor3b_wx109 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps110 = multm_reduce_mulb0_add3b_xor3b_wx110 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps111 = multm_reduce_mulb0_sq112 ^ multm_reduce_mulb0_cq111;
  assign multm_reduce_mulb0_ps112 = multm_reduce_mulb0_sq113 ^ multm_reduce_mulb0_cq112;
  assign multm_reduce_mulb0_ps113 = multm_reduce_mulb0_sq114 ^ multm_reduce_mulb0_cq113;
  assign multm_reduce_mulb0_ps114 = multm_reduce_mulb0_add3b_xor3b_wx114 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps115 = multm_reduce_mulb0_sq116 ^ multm_reduce_mulb0_cq115;
  assign multm_reduce_mulb0_ps116 = multm_reduce_mulb0_sq117 ^ multm_reduce_mulb0_cq116;
  assign multm_reduce_mulb0_ps117 = multm_reduce_mulb0_add3b_xor3b_wx117 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps118 = multm_reduce_mulb0_add3b_xor3b_wx118 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps119 = multm_reduce_mulb0_sq120 ^ multm_reduce_mulb0_cq119;
  assign multm_reduce_mulb0_ps120 = multm_reduce_mulb0_add3b_xor3b_wx120 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps121 = multm_reduce_mulb0_sq122 ^ multm_reduce_mulb0_cq121;
  assign multm_reduce_mulb0_ps122 = multm_reduce_mulb0_add3b_xor3b_wx122 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps123 = multm_reduce_mulb0_add3b_xor3b_wx123 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps124 = multm_reduce_mulb0_sq125 ^ multm_reduce_mulb0_cq124;
  assign multm_reduce_mulb0_ps125 = multm_reduce_mulb0_sq126 ^ multm_reduce_mulb0_cq125;
  assign multm_reduce_mulb0_ps126 = multm_reduce_mulb0_sq127 ^ multm_reduce_mulb0_cq126;
  assign multm_reduce_mulb0_ps127 = multm_reduce_mulb0_add3b_xor3b_wx127 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps128 = multm_reduce_mulb0_add3b_xor3b_wx128 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps129 = multm_reduce_mulb0_sq130 ^ multm_reduce_mulb0_cq129;
  assign multm_reduce_mulb0_ps130 = multm_reduce_mulb0_sq131 ^ multm_reduce_mulb0_cq130;
  assign multm_reduce_mulb0_ps131 = multm_reduce_mulb0_add3b_xor3b_wx131 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps132 = multm_reduce_mulb0_sq133 ^ multm_reduce_mulb0_cq132;
  assign multm_reduce_mulb0_ps133 = multm_reduce_mulb0_sq134 ^ multm_reduce_mulb0_cq133;
  assign multm_reduce_mulb0_ps134 = multm_reduce_mulb0_add3b_xor3b_wx134 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps135 = multm_reduce_mulb0_add3b_xor3b_wx135 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps136 = multm_reduce_mulb0_add3b_xor3b_wx136 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps137 = multm_reduce_mulb0_sq138 ^ multm_reduce_mulb0_cq137;
  assign multm_reduce_mulb0_ps138 = multm_reduce_mulb0_add3b_xor3b_wx138 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps139 = multm_reduce_mulb0_sq140 ^ multm_reduce_mulb0_cq139;
  assign multm_reduce_mulb0_ps140 = multm_reduce_mulb0_add3b_xor3b_wx140 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps141 = multm_reduce_mulb0_sq142 ^ multm_reduce_mulb0_cq141;
  assign multm_reduce_mulb0_ps142 = multm_reduce_mulb0_sq143 ^ multm_reduce_mulb0_cq142;
  assign multm_reduce_mulb0_ps143 = multm_reduce_mulb0_sq144 ^ multm_reduce_mulb0_cq143;
  assign multm_reduce_mulb0_ps144 = multm_reduce_mulb0_sq145 ^ multm_reduce_mulb0_cq144;
  assign multm_reduce_mulb0_ps145 = multm_reduce_mulb0_sq146 ^ multm_reduce_mulb0_cq145;
  assign multm_reduce_mulb0_ps146 = multm_reduce_mulb0_add3b_xor3b_wx146 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps147 = multm_reduce_mulb0_add3b_xor3b_wx147 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps148 = multm_reduce_mulb0_add3b_xor3b_wx148 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps149 = multm_reduce_mulb0_add3b_xor3b_wx149 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps150 = multm_reduce_mulb0_sq151 ^ multm_reduce_mulb0_cq150;
  assign multm_reduce_mulb0_ps151 = multm_reduce_mulb0_sq152 ^ multm_reduce_mulb0_cq151;
  assign multm_reduce_mulb0_ps152 = multm_reduce_mulb0_add3b_xor3b_wx152 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps153 = multm_reduce_mulb0_add3b_xor3b_wx153 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps154 = multm_reduce_mulb0_sq155 ^ multm_reduce_mulb0_cq154;
  assign multm_reduce_mulb0_ps155 = multm_reduce_mulb0_sq156 ^ multm_reduce_mulb0_cq155;
  assign multm_reduce_mulb0_ps156 = multm_reduce_mulb0_add3b_xor3b_wx156 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps157 = multm_reduce_mulb0_add3b_xor3b_wx157 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps158 = multm_reduce_mulb0_add3b_xor3b_wx158 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps159 = multm_reduce_mulb0_add3b_xor3b_wx159 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps160 = multm_reduce_mulb0_add3b_xor3b_wx160 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps161 = multm_reduce_mulb0_sq162 ^ multm_reduce_mulb0_cq161;
  assign multm_reduce_mulb0_ps162 = multm_reduce_mulb0_add3b_xor3b_wx162 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps163 = multm_reduce_mulb0_add3b_xor3b_wx163 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps164 = multm_reduce_mulb0_sq165 ^ multm_reduce_mulb0_cq164;
  assign multm_reduce_mulb0_ps165 = multm_reduce_mulb0_sq166 ^ multm_reduce_mulb0_cq165;
  assign multm_reduce_mulb0_ps166 = multm_reduce_mulb0_sq167 ^ multm_reduce_mulb0_cq166;
  assign multm_reduce_mulb0_ps167 = multm_reduce_mulb0_sq168 ^ multm_reduce_mulb0_cq167;
  assign multm_reduce_mulb0_ps168 = multm_reduce_mulb0_add3b_xor3b_wx168 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps169 = multm_reduce_mulb0_sq170 ^ multm_reduce_mulb0_cq169;
  assign multm_reduce_mulb0_ps170 = multm_reduce_mulb0_add3b_xor3b_wx170 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps171 = multm_reduce_mulb0_add3b_xor3b_wx171 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps172 = multm_reduce_mulb0_add3b_xor3b_wx172 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps173 = multm_reduce_mulb0_add3b_xor3b_wx173 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps174 = multm_reduce_mulb0_sq175 ^ multm_reduce_mulb0_cq174;
  assign multm_reduce_mulb0_ps175 = multm_reduce_mulb0_add3b_xor3b_wx175 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps176 = multm_reduce_mulb0_sq177 ^ multm_reduce_mulb0_cq176;
  assign multm_reduce_mulb0_ps177 = multm_reduce_mulb0_add3b_xor3b_wx177 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps178 = multm_reduce_mulb0_add3b_xor3b_wx178 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps179 = multm_reduce_mulb0_sq180 ^ multm_reduce_mulb0_cq179;
  assign multm_reduce_mulb0_ps180 = multm_reduce_mulb0_sq181 ^ multm_reduce_mulb0_cq180;
  assign multm_reduce_mulb0_ps181 = multm_reduce_mulb0_add3b_xor3b_wx181 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps182 = multm_reduce_mulb0_add3b_xor3b_wx182 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_ps183 = multm_reduce_mulb0_add3b_xor3b_wx183 ^ multm_reduce_sa5;
  assign multm_reduce_mulb0_sq0 = xn1 & multm_reduce_mulb0_sp0;
  assign multm_reduce_mulb0_sq1 = xn1 & multm_reduce_mulb0_sp1;
  assign multm_reduce_mulb0_sq2 = xn1 & multm_reduce_mulb0_sp2;
  assign multm_reduce_mulb0_sq3 = xn1 & multm_reduce_mulb0_sp3;
  assign multm_reduce_mulb0_sq4 = xn1 & multm_reduce_mulb0_sp4;
  assign multm_reduce_mulb0_sq5 = xn1 & multm_reduce_mulb0_sp5;
  assign multm_reduce_mulb0_sq6 = xn1 & multm_reduce_mulb0_sp6;
  assign multm_reduce_mulb0_sq7 = xn1 & multm_reduce_mulb0_sp7;
  assign multm_reduce_mulb0_sq8 = xn1 & multm_reduce_mulb0_sp8;
  assign multm_reduce_mulb0_sq9 = xn1 & multm_reduce_mulb0_sp9;
  assign multm_reduce_mulb0_sq10 = xn1 & multm_reduce_mulb0_sp10;
  assign multm_reduce_mulb0_sq11 = xn1 & multm_reduce_mulb0_sp11;
  assign multm_reduce_mulb0_sq12 = xn1 & multm_reduce_mulb0_sp12;
  assign multm_reduce_mulb0_sq13 = xn1 & multm_reduce_mulb0_sp13;
  assign multm_reduce_mulb0_sq14 = xn1 & multm_reduce_mulb0_sp14;
  assign multm_reduce_mulb0_sq15 = xn1 & multm_reduce_mulb0_sp15;
  assign multm_reduce_mulb0_sq16 = xn1 & multm_reduce_mulb0_sp16;
  assign multm_reduce_mulb0_sq17 = xn1 & multm_reduce_mulb0_sp17;
  assign multm_reduce_mulb0_sq18 = xn1 & multm_reduce_mulb0_sp18;
  assign multm_reduce_mulb0_sq19 = xn1 & multm_reduce_mulb0_sp19;
  assign multm_reduce_mulb0_sq20 = xn1 & multm_reduce_mulb0_sp20;
  assign multm_reduce_mulb0_sq21 = xn1 & multm_reduce_mulb0_sp21;
  assign multm_reduce_mulb0_sq22 = xn1 & multm_reduce_mulb0_sp22;
  assign multm_reduce_mulb0_sq23 = xn1 & multm_reduce_mulb0_sp23;
  assign multm_reduce_mulb0_sq24 = xn1 & multm_reduce_mulb0_sp24;
  assign multm_reduce_mulb0_sq25 = xn1 & multm_reduce_mulb0_sp25;
  assign multm_reduce_mulb0_sq26 = xn1 & multm_reduce_mulb0_sp26;
  assign multm_reduce_mulb0_sq27 = xn1 & multm_reduce_mulb0_sp27;
  assign multm_reduce_mulb0_sq28 = xn1 & multm_reduce_mulb0_sp28;
  assign multm_reduce_mulb0_sq29 = xn1 & multm_reduce_mulb0_sp29;
  assign multm_reduce_mulb0_sq30 = xn1 & multm_reduce_mulb0_sp30;
  assign multm_reduce_mulb0_sq31 = xn1 & multm_reduce_mulb0_sp31;
  assign multm_reduce_mulb0_sq32 = xn1 & multm_reduce_mulb0_sp32;
  assign multm_reduce_mulb0_sq33 = xn1 & multm_reduce_mulb0_sp33;
  assign multm_reduce_mulb0_sq34 = xn1 & multm_reduce_mulb0_sp34;
  assign multm_reduce_mulb0_sq35 = xn1 & multm_reduce_mulb0_sp35;
  assign multm_reduce_mulb0_sq36 = xn1 & multm_reduce_mulb0_sp36;
  assign multm_reduce_mulb0_sq37 = xn1 & multm_reduce_mulb0_sp37;
  assign multm_reduce_mulb0_sq38 = xn1 & multm_reduce_mulb0_sp38;
  assign multm_reduce_mulb0_sq39 = xn1 & multm_reduce_mulb0_sp39;
  assign multm_reduce_mulb0_sq40 = xn1 & multm_reduce_mulb0_sp40;
  assign multm_reduce_mulb0_sq41 = xn1 & multm_reduce_mulb0_sp41;
  assign multm_reduce_mulb0_sq42 = xn1 & multm_reduce_mulb0_sp42;
  assign multm_reduce_mulb0_sq43 = xn1 & multm_reduce_mulb0_sp43;
  assign multm_reduce_mulb0_sq44 = xn1 & multm_reduce_mulb0_sp44;
  assign multm_reduce_mulb0_sq45 = xn1 & multm_reduce_mulb0_sp45;
  assign multm_reduce_mulb0_sq46 = xn1 & multm_reduce_mulb0_sp46;
  assign multm_reduce_mulb0_sq47 = xn1 & multm_reduce_mulb0_sp47;
  assign multm_reduce_mulb0_sq48 = xn1 & multm_reduce_mulb0_sp48;
  assign multm_reduce_mulb0_sq49 = xn1 & multm_reduce_mulb0_sp49;
  assign multm_reduce_mulb0_sq50 = xn1 & multm_reduce_mulb0_sp50;
  assign multm_reduce_mulb0_sq51 = xn1 & multm_reduce_mulb0_sp51;
  assign multm_reduce_mulb0_sq52 = xn1 & multm_reduce_mulb0_sp52;
  assign multm_reduce_mulb0_sq53 = xn1 & multm_reduce_mulb0_sp53;
  assign multm_reduce_mulb0_sq54 = xn1 & multm_reduce_mulb0_sp54;
  assign multm_reduce_mulb0_sq55 = xn1 & multm_reduce_mulb0_sp55;
  assign multm_reduce_mulb0_sq56 = xn1 & multm_reduce_mulb0_sp56;
  assign multm_reduce_mulb0_sq57 = xn1 & multm_reduce_mulb0_sp57;
  assign multm_reduce_mulb0_sq58 = xn1 & multm_reduce_mulb0_sp58;
  assign multm_reduce_mulb0_sq59 = xn1 & multm_reduce_mulb0_sp59;
  assign multm_reduce_mulb0_sq60 = xn1 & multm_reduce_mulb0_sp60;
  assign multm_reduce_mulb0_sq61 = xn1 & multm_reduce_mulb0_sp61;
  assign multm_reduce_mulb0_sq62 = xn1 & multm_reduce_mulb0_sp62;
  assign multm_reduce_mulb0_sq63 = xn1 & multm_reduce_mulb0_sp63;
  assign multm_reduce_mulb0_sq64 = xn1 & multm_reduce_mulb0_sp64;
  assign multm_reduce_mulb0_sq65 = xn1 & multm_reduce_mulb0_sp65;
  assign multm_reduce_mulb0_sq66 = xn1 & multm_reduce_mulb0_sp66;
  assign multm_reduce_mulb0_sq67 = xn1 & multm_reduce_mulb0_sp67;
  assign multm_reduce_mulb0_sq68 = xn1 & multm_reduce_mulb0_sp68;
  assign multm_reduce_mulb0_sq69 = xn1 & multm_reduce_mulb0_sp69;
  assign multm_reduce_mulb0_sq70 = xn1 & multm_reduce_mulb0_sp70;
  assign multm_reduce_mulb0_sq71 = xn1 & multm_reduce_mulb0_sp71;
  assign multm_reduce_mulb0_sq72 = xn1 & multm_reduce_mulb0_sp72;
  assign multm_reduce_mulb0_sq73 = xn1 & multm_reduce_mulb0_sp73;
  assign multm_reduce_mulb0_sq74 = xn1 & multm_reduce_mulb0_sp74;
  assign multm_reduce_mulb0_sq75 = xn1 & multm_reduce_mulb0_sp75;
  assign multm_reduce_mulb0_sq76 = xn1 & multm_reduce_mulb0_sp76;
  assign multm_reduce_mulb0_sq77 = xn1 & multm_reduce_mulb0_sp77;
  assign multm_reduce_mulb0_sq78 = xn1 & multm_reduce_mulb0_sp78;
  assign multm_reduce_mulb0_sq79 = xn1 & multm_reduce_mulb0_sp79;
  assign multm_reduce_mulb0_sq80 = xn1 & multm_reduce_mulb0_sp80;
  assign multm_reduce_mulb0_sq81 = xn1 & multm_reduce_mulb0_sp81;
  assign multm_reduce_mulb0_sq82 = xn1 & multm_reduce_mulb0_sp82;
  assign multm_reduce_mulb0_sq83 = xn1 & multm_reduce_mulb0_sp83;
  assign multm_reduce_mulb0_sq84 = xn1 & multm_reduce_mulb0_sp84;
  assign multm_reduce_mulb0_sq85 = xn1 & multm_reduce_mulb0_sp85;
  assign multm_reduce_mulb0_sq86 = xn1 & multm_reduce_mulb0_sp86;
  assign multm_reduce_mulb0_sq87 = xn1 & multm_reduce_mulb0_sp87;
  assign multm_reduce_mulb0_sq88 = xn1 & multm_reduce_mulb0_sp88;
  assign multm_reduce_mulb0_sq89 = xn1 & multm_reduce_mulb0_sp89;
  assign multm_reduce_mulb0_sq90 = xn1 & multm_reduce_mulb0_sp90;
  assign multm_reduce_mulb0_sq91 = xn1 & multm_reduce_mulb0_sp91;
  assign multm_reduce_mulb0_sq92 = xn1 & multm_reduce_mulb0_sp92;
  assign multm_reduce_mulb0_sq93 = xn1 & multm_reduce_mulb0_sp93;
  assign multm_reduce_mulb0_sq94 = xn1 & multm_reduce_mulb0_sp94;
  assign multm_reduce_mulb0_sq95 = xn1 & multm_reduce_mulb0_sp95;
  assign multm_reduce_mulb0_sq96 = xn1 & multm_reduce_mulb0_sp96;
  assign multm_reduce_mulb0_sq97 = xn1 & multm_reduce_mulb0_sp97;
  assign multm_reduce_mulb0_sq98 = xn1 & multm_reduce_mulb0_sp98;
  assign multm_reduce_mulb0_sq99 = xn1 & multm_reduce_mulb0_sp99;
  assign multm_reduce_mulb0_sq100 = xn1 & multm_reduce_mulb0_sp100;
  assign multm_reduce_mulb0_sq101 = xn1 & multm_reduce_mulb0_sp101;
  assign multm_reduce_mulb0_sq102 = xn1 & multm_reduce_mulb0_sp102;
  assign multm_reduce_mulb0_sq103 = xn1 & multm_reduce_mulb0_sp103;
  assign multm_reduce_mulb0_sq104 = xn1 & multm_reduce_mulb0_sp104;
  assign multm_reduce_mulb0_sq105 = xn1 & multm_reduce_mulb0_sp105;
  assign multm_reduce_mulb0_sq106 = xn1 & multm_reduce_mulb0_sp106;
  assign multm_reduce_mulb0_sq107 = xn1 & multm_reduce_mulb0_sp107;
  assign multm_reduce_mulb0_sq108 = xn1 & multm_reduce_mulb0_sp108;
  assign multm_reduce_mulb0_sq109 = xn1 & multm_reduce_mulb0_sp109;
  assign multm_reduce_mulb0_sq110 = xn1 & multm_reduce_mulb0_sp110;
  assign multm_reduce_mulb0_sq111 = xn1 & multm_reduce_mulb0_sp111;
  assign multm_reduce_mulb0_sq112 = xn1 & multm_reduce_mulb0_sp112;
  assign multm_reduce_mulb0_sq113 = xn1 & multm_reduce_mulb0_sp113;
  assign multm_reduce_mulb0_sq114 = xn1 & multm_reduce_mulb0_sp114;
  assign multm_reduce_mulb0_sq115 = xn1 & multm_reduce_mulb0_sp115;
  assign multm_reduce_mulb0_sq116 = xn1 & multm_reduce_mulb0_sp116;
  assign multm_reduce_mulb0_sq117 = xn1 & multm_reduce_mulb0_sp117;
  assign multm_reduce_mulb0_sq118 = xn1 & multm_reduce_mulb0_sp118;
  assign multm_reduce_mulb0_sq119 = xn1 & multm_reduce_mulb0_sp119;
  assign multm_reduce_mulb0_sq120 = xn1 & multm_reduce_mulb0_sp120;
  assign multm_reduce_mulb0_sq121 = xn1 & multm_reduce_mulb0_sp121;
  assign multm_reduce_mulb0_sq122 = xn1 & multm_reduce_mulb0_sp122;
  assign multm_reduce_mulb0_sq123 = xn1 & multm_reduce_mulb0_sp123;
  assign multm_reduce_mulb0_sq124 = xn1 & multm_reduce_mulb0_sp124;
  assign multm_reduce_mulb0_sq125 = xn1 & multm_reduce_mulb0_sp125;
  assign multm_reduce_mulb0_sq126 = xn1 & multm_reduce_mulb0_sp126;
  assign multm_reduce_mulb0_sq127 = xn1 & multm_reduce_mulb0_sp127;
  assign multm_reduce_mulb0_sq128 = xn1 & multm_reduce_mulb0_sp128;
  assign multm_reduce_mulb0_sq129 = xn1 & multm_reduce_mulb0_sp129;
  assign multm_reduce_mulb0_sq130 = xn1 & multm_reduce_mulb0_sp130;
  assign multm_reduce_mulb0_sq131 = xn1 & multm_reduce_mulb0_sp131;
  assign multm_reduce_mulb0_sq132 = xn1 & multm_reduce_mulb0_sp132;
  assign multm_reduce_mulb0_sq133 = xn1 & multm_reduce_mulb0_sp133;
  assign multm_reduce_mulb0_sq134 = xn1 & multm_reduce_mulb0_sp134;
  assign multm_reduce_mulb0_sq135 = xn1 & multm_reduce_mulb0_sp135;
  assign multm_reduce_mulb0_sq136 = xn1 & multm_reduce_mulb0_sp136;
  assign multm_reduce_mulb0_sq137 = xn1 & multm_reduce_mulb0_sp137;
  assign multm_reduce_mulb0_sq138 = xn1 & multm_reduce_mulb0_sp138;
  assign multm_reduce_mulb0_sq139 = xn1 & multm_reduce_mulb0_sp139;
  assign multm_reduce_mulb0_sq140 = xn1 & multm_reduce_mulb0_sp140;
  assign multm_reduce_mulb0_sq141 = xn1 & multm_reduce_mulb0_sp141;
  assign multm_reduce_mulb0_sq142 = xn1 & multm_reduce_mulb0_sp142;
  assign multm_reduce_mulb0_sq143 = xn1 & multm_reduce_mulb0_sp143;
  assign multm_reduce_mulb0_sq144 = xn1 & multm_reduce_mulb0_sp144;
  assign multm_reduce_mulb0_sq145 = xn1 & multm_reduce_mulb0_sp145;
  assign multm_reduce_mulb0_sq146 = xn1 & multm_reduce_mulb0_sp146;
  assign multm_reduce_mulb0_sq147 = xn1 & multm_reduce_mulb0_sp147;
  assign multm_reduce_mulb0_sq148 = xn1 & multm_reduce_mulb0_sp148;
  assign multm_reduce_mulb0_sq149 = xn1 & multm_reduce_mulb0_sp149;
  assign multm_reduce_mulb0_sq150 = xn1 & multm_reduce_mulb0_sp150;
  assign multm_reduce_mulb0_sq151 = xn1 & multm_reduce_mulb0_sp151;
  assign multm_reduce_mulb0_sq152 = xn1 & multm_reduce_mulb0_sp152;
  assign multm_reduce_mulb0_sq153 = xn1 & multm_reduce_mulb0_sp153;
  assign multm_reduce_mulb0_sq154 = xn1 & multm_reduce_mulb0_sp154;
  assign multm_reduce_mulb0_sq155 = xn1 & multm_reduce_mulb0_sp155;
  assign multm_reduce_mulb0_sq156 = xn1 & multm_reduce_mulb0_sp156;
  assign multm_reduce_mulb0_sq157 = xn1 & multm_reduce_mulb0_sp157;
  assign multm_reduce_mulb0_sq158 = xn1 & multm_reduce_mulb0_sp158;
  assign multm_reduce_mulb0_sq159 = xn1 & multm_reduce_mulb0_sp159;
  assign multm_reduce_mulb0_sq160 = xn1 & multm_reduce_mulb0_sp160;
  assign multm_reduce_mulb0_sq161 = xn1 & multm_reduce_mulb0_sp161;
  assign multm_reduce_mulb0_sq162 = xn1 & multm_reduce_mulb0_sp162;
  assign multm_reduce_mulb0_sq163 = xn1 & multm_reduce_mulb0_sp163;
  assign multm_reduce_mulb0_sq164 = xn1 & multm_reduce_mulb0_sp164;
  assign multm_reduce_mulb0_sq165 = xn1 & multm_reduce_mulb0_sp165;
  assign multm_reduce_mulb0_sq166 = xn1 & multm_reduce_mulb0_sp166;
  assign multm_reduce_mulb0_sq167 = xn1 & multm_reduce_mulb0_sp167;
  assign multm_reduce_mulb0_sq168 = xn1 & multm_reduce_mulb0_sp168;
  assign multm_reduce_mulb0_sq169 = xn1 & multm_reduce_mulb0_sp169;
  assign multm_reduce_mulb0_sq170 = xn1 & multm_reduce_mulb0_sp170;
  assign multm_reduce_mulb0_sq171 = xn1 & multm_reduce_mulb0_sp171;
  assign multm_reduce_mulb0_sq172 = xn1 & multm_reduce_mulb0_sp172;
  assign multm_reduce_mulb0_sq173 = xn1 & multm_reduce_mulb0_sp173;
  assign multm_reduce_mulb0_sq174 = xn1 & multm_reduce_mulb0_sp174;
  assign multm_reduce_mulb0_sq175 = xn1 & multm_reduce_mulb0_sp175;
  assign multm_reduce_mulb0_sq176 = xn1 & multm_reduce_mulb0_sp176;
  assign multm_reduce_mulb0_sq177 = xn1 & multm_reduce_mulb0_sp177;
  assign multm_reduce_mulb0_sq178 = xn1 & multm_reduce_mulb0_sp178;
  assign multm_reduce_mulb0_sq179 = xn1 & multm_reduce_mulb0_sp179;
  assign multm_reduce_mulb0_sq180 = xn1 & multm_reduce_mulb0_sp180;
  assign multm_reduce_mulb0_sq181 = xn1 & multm_reduce_mulb0_sp181;
  assign multm_reduce_mulb0_sq182 = xn1 & multm_reduce_mulb0_sp182;
  assign multm_reduce_mulb0_sq183 = xn1 & multm_reduce_mulb0_sp183;
  assign multm_reduce_mulb0_sq184 = xn1 & multm_reduce_mulb0_sp184;
  assign multm_reduce_mulb1_add3_maj3_or3_wx = multm_reduce_mulb1_add3_maj3_wx | multm_reduce_mulb1_add3_maj3_wy;
  assign multm_reduce_mulb1_add3_maj3_wx = multm_reduce_qb2 & multm_reduce_mulb1_cq182;
  assign multm_reduce_mulb1_add3_maj3_wy = multm_reduce_qb2 & multm_reduce_mulb1_pc182;
  assign multm_reduce_mulb1_add3_maj3_xy = multm_reduce_mulb1_cq182 & multm_reduce_mulb1_pc182;
  assign multm_reduce_mulb1_add3_xor3_wx = multm_reduce_qb2 ^ multm_reduce_mulb1_cq182;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx0 = multm_reduce_mulb1_add3b_maj3b_wx0 | multm_reduce_mulb1_add3b_maj3b_wy0;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx1 = multm_reduce_mulb1_add3b_maj3b_wx1 | multm_reduce_mulb1_add3b_maj3b_wy1;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx4 = multm_reduce_mulb1_add3b_maj3b_wx4 | multm_reduce_mulb1_add3b_maj3b_wy4;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx5 = multm_reduce_mulb1_add3b_maj3b_wx5 | multm_reduce_mulb1_add3b_maj3b_wy5;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx6 = multm_reduce_mulb1_add3b_maj3b_wx6 | multm_reduce_mulb1_add3b_maj3b_wy6;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx7 = multm_reduce_mulb1_add3b_maj3b_wx7 | multm_reduce_mulb1_add3b_maj3b_wy7;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx10 = multm_reduce_mulb1_add3b_maj3b_wx10 | multm_reduce_mulb1_add3b_maj3b_wy10;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx12 = multm_reduce_mulb1_add3b_maj3b_wx12 | multm_reduce_mulb1_add3b_maj3b_wy12;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx18 = multm_reduce_mulb1_add3b_maj3b_wx18 | multm_reduce_mulb1_add3b_maj3b_wy18;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx20 = multm_reduce_mulb1_add3b_maj3b_wx20 | multm_reduce_mulb1_add3b_maj3b_wy20;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx22 = multm_reduce_mulb1_add3b_maj3b_wx22 | multm_reduce_mulb1_add3b_maj3b_wy22;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx23 = multm_reduce_mulb1_add3b_maj3b_wx23 | multm_reduce_mulb1_add3b_maj3b_wy23;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx24 = multm_reduce_mulb1_add3b_maj3b_wx24 | multm_reduce_mulb1_add3b_maj3b_wy24;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx28 = multm_reduce_mulb1_add3b_maj3b_wx28 | multm_reduce_mulb1_add3b_maj3b_wy28;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx30 = multm_reduce_mulb1_add3b_maj3b_wx30 | multm_reduce_mulb1_add3b_maj3b_wy30;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx32 = multm_reduce_mulb1_add3b_maj3b_wx32 | multm_reduce_mulb1_add3b_maj3b_wy32;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx34 = multm_reduce_mulb1_add3b_maj3b_wx34 | multm_reduce_mulb1_add3b_maj3b_wy34;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx37 = multm_reduce_mulb1_add3b_maj3b_wx37 | multm_reduce_mulb1_add3b_maj3b_wy37;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx40 = multm_reduce_mulb1_add3b_maj3b_wx40 | multm_reduce_mulb1_add3b_maj3b_wy40;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx41 = multm_reduce_mulb1_add3b_maj3b_wx41 | multm_reduce_mulb1_add3b_maj3b_wy41;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx42 = multm_reduce_mulb1_add3b_maj3b_wx42 | multm_reduce_mulb1_add3b_maj3b_wy42;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx43 = multm_reduce_mulb1_add3b_maj3b_wx43 | multm_reduce_mulb1_add3b_maj3b_wy43;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx47 = multm_reduce_mulb1_add3b_maj3b_wx47 | multm_reduce_mulb1_add3b_maj3b_wy47;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx48 = multm_reduce_mulb1_add3b_maj3b_wx48 | multm_reduce_mulb1_add3b_maj3b_wy48;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx51 = multm_reduce_mulb1_add3b_maj3b_wx51 | multm_reduce_mulb1_add3b_maj3b_wy51;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx52 = multm_reduce_mulb1_add3b_maj3b_wx52 | multm_reduce_mulb1_add3b_maj3b_wy52;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx53 = multm_reduce_mulb1_add3b_maj3b_wx53 | multm_reduce_mulb1_add3b_maj3b_wy53;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx54 = multm_reduce_mulb1_add3b_maj3b_wx54 | multm_reduce_mulb1_add3b_maj3b_wy54;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx55 = multm_reduce_mulb1_add3b_maj3b_wx55 | multm_reduce_mulb1_add3b_maj3b_wy55;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx57 = multm_reduce_mulb1_add3b_maj3b_wx57 | multm_reduce_mulb1_add3b_maj3b_wy57;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx62 = multm_reduce_mulb1_add3b_maj3b_wx62 | multm_reduce_mulb1_add3b_maj3b_wy62;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx66 = multm_reduce_mulb1_add3b_maj3b_wx66 | multm_reduce_mulb1_add3b_maj3b_wy66;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx68 = multm_reduce_mulb1_add3b_maj3b_wx68 | multm_reduce_mulb1_add3b_maj3b_wy68;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx69 = multm_reduce_mulb1_add3b_maj3b_wx69 | multm_reduce_mulb1_add3b_maj3b_wy69;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx71 = multm_reduce_mulb1_add3b_maj3b_wx71 | multm_reduce_mulb1_add3b_maj3b_wy71;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx73 = multm_reduce_mulb1_add3b_maj3b_wx73 | multm_reduce_mulb1_add3b_maj3b_wy73;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx74 = multm_reduce_mulb1_add3b_maj3b_wx74 | multm_reduce_mulb1_add3b_maj3b_wy74;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx79 = multm_reduce_mulb1_add3b_maj3b_wx79 | multm_reduce_mulb1_add3b_maj3b_wy79;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx80 = multm_reduce_mulb1_add3b_maj3b_wx80 | multm_reduce_mulb1_add3b_maj3b_wy80;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx82 = multm_reduce_mulb1_add3b_maj3b_wx82 | multm_reduce_mulb1_add3b_maj3b_wy82;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx86 = multm_reduce_mulb1_add3b_maj3b_wx86 | multm_reduce_mulb1_add3b_maj3b_wy86;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx88 = multm_reduce_mulb1_add3b_maj3b_wx88 | multm_reduce_mulb1_add3b_maj3b_wy88;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx90 = multm_reduce_mulb1_add3b_maj3b_wx90 | multm_reduce_mulb1_add3b_maj3b_wy90;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx91 = multm_reduce_mulb1_add3b_maj3b_wx91 | multm_reduce_mulb1_add3b_maj3b_wy91;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx96 = multm_reduce_mulb1_add3b_maj3b_wx96 | multm_reduce_mulb1_add3b_maj3b_wy96;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx99 = multm_reduce_mulb1_add3b_maj3b_wx99 | multm_reduce_mulb1_add3b_maj3b_wy99;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx100 = multm_reduce_mulb1_add3b_maj3b_wx100 | multm_reduce_mulb1_add3b_maj3b_wy100;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx101 = multm_reduce_mulb1_add3b_maj3b_wx101 | multm_reduce_mulb1_add3b_maj3b_wy101;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx102 = multm_reduce_mulb1_add3b_maj3b_wx102 | multm_reduce_mulb1_add3b_maj3b_wy102;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx104 = multm_reduce_mulb1_add3b_maj3b_wx104 | multm_reduce_mulb1_add3b_maj3b_wy104;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx105 = multm_reduce_mulb1_add3b_maj3b_wx105 | multm_reduce_mulb1_add3b_maj3b_wy105;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx107 = multm_reduce_mulb1_add3b_maj3b_wx107 | multm_reduce_mulb1_add3b_maj3b_wy107;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx108 = multm_reduce_mulb1_add3b_maj3b_wx108 | multm_reduce_mulb1_add3b_maj3b_wy108;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx109 = multm_reduce_mulb1_add3b_maj3b_wx109 | multm_reduce_mulb1_add3b_maj3b_wy109;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx110 = multm_reduce_mulb1_add3b_maj3b_wx110 | multm_reduce_mulb1_add3b_maj3b_wy110;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx112 = multm_reduce_mulb1_add3b_maj3b_wx112 | multm_reduce_mulb1_add3b_maj3b_wy112;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx114 = multm_reduce_mulb1_add3b_maj3b_wx114 | multm_reduce_mulb1_add3b_maj3b_wy114;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx117 = multm_reduce_mulb1_add3b_maj3b_wx117 | multm_reduce_mulb1_add3b_maj3b_wy117;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx118 = multm_reduce_mulb1_add3b_maj3b_wx118 | multm_reduce_mulb1_add3b_maj3b_wy118;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx119 = multm_reduce_mulb1_add3b_maj3b_wx119 | multm_reduce_mulb1_add3b_maj3b_wy119;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx120 = multm_reduce_mulb1_add3b_maj3b_wx120 | multm_reduce_mulb1_add3b_maj3b_wy120;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx121 = multm_reduce_mulb1_add3b_maj3b_wx121 | multm_reduce_mulb1_add3b_maj3b_wy121;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx122 = multm_reduce_mulb1_add3b_maj3b_wx122 | multm_reduce_mulb1_add3b_maj3b_wy122;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx123 = multm_reduce_mulb1_add3b_maj3b_wx123 | multm_reduce_mulb1_add3b_maj3b_wy123;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx128 = multm_reduce_mulb1_add3b_maj3b_wx128 | multm_reduce_mulb1_add3b_maj3b_wy128;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx130 = multm_reduce_mulb1_add3b_maj3b_wx130 | multm_reduce_mulb1_add3b_maj3b_wy130;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx132 = multm_reduce_mulb1_add3b_maj3b_wx132 | multm_reduce_mulb1_add3b_maj3b_wy132;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx135 = multm_reduce_mulb1_add3b_maj3b_wx135 | multm_reduce_mulb1_add3b_maj3b_wy135;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx136 = multm_reduce_mulb1_add3b_maj3b_wx136 | multm_reduce_mulb1_add3b_maj3b_wy136;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx140 = multm_reduce_mulb1_add3b_maj3b_wx140 | multm_reduce_mulb1_add3b_maj3b_wy140;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx141 = multm_reduce_mulb1_add3b_maj3b_wx141 | multm_reduce_mulb1_add3b_maj3b_wy141;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx142 = multm_reduce_mulb1_add3b_maj3b_wx142 | multm_reduce_mulb1_add3b_maj3b_wy142;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx143 = multm_reduce_mulb1_add3b_maj3b_wx143 | multm_reduce_mulb1_add3b_maj3b_wy143;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx144 = multm_reduce_mulb1_add3b_maj3b_wx144 | multm_reduce_mulb1_add3b_maj3b_wy144;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx147 = multm_reduce_mulb1_add3b_maj3b_wx147 | multm_reduce_mulb1_add3b_maj3b_wy147;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx150 = multm_reduce_mulb1_add3b_maj3b_wx150 | multm_reduce_mulb1_add3b_maj3b_wy150;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx151 = multm_reduce_mulb1_add3b_maj3b_wx151 | multm_reduce_mulb1_add3b_maj3b_wy151;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx152 = multm_reduce_mulb1_add3b_maj3b_wx152 | multm_reduce_mulb1_add3b_maj3b_wy152;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx153 = multm_reduce_mulb1_add3b_maj3b_wx153 | multm_reduce_mulb1_add3b_maj3b_wy153;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx155 = multm_reduce_mulb1_add3b_maj3b_wx155 | multm_reduce_mulb1_add3b_maj3b_wy155;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx156 = multm_reduce_mulb1_add3b_maj3b_wx156 | multm_reduce_mulb1_add3b_maj3b_wy156;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx157 = multm_reduce_mulb1_add3b_maj3b_wx157 | multm_reduce_mulb1_add3b_maj3b_wy157;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx158 = multm_reduce_mulb1_add3b_maj3b_wx158 | multm_reduce_mulb1_add3b_maj3b_wy158;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx159 = multm_reduce_mulb1_add3b_maj3b_wx159 | multm_reduce_mulb1_add3b_maj3b_wy159;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx160 = multm_reduce_mulb1_add3b_maj3b_wx160 | multm_reduce_mulb1_add3b_maj3b_wy160;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx162 = multm_reduce_mulb1_add3b_maj3b_wx162 | multm_reduce_mulb1_add3b_maj3b_wy162;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx166 = multm_reduce_mulb1_add3b_maj3b_wx166 | multm_reduce_mulb1_add3b_maj3b_wy166;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx171 = multm_reduce_mulb1_add3b_maj3b_wx171 | multm_reduce_mulb1_add3b_maj3b_wy171;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx172 = multm_reduce_mulb1_add3b_maj3b_wx172 | multm_reduce_mulb1_add3b_maj3b_wy172;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx173 = multm_reduce_mulb1_add3b_maj3b_wx173 | multm_reduce_mulb1_add3b_maj3b_wy173;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx174 = multm_reduce_mulb1_add3b_maj3b_wx174 | multm_reduce_mulb1_add3b_maj3b_wy174;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx175 = multm_reduce_mulb1_add3b_maj3b_wx175 | multm_reduce_mulb1_add3b_maj3b_wy175;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx179 = multm_reduce_mulb1_add3b_maj3b_wx179 | multm_reduce_mulb1_add3b_maj3b_wy179;
  assign multm_reduce_mulb1_add3b_maj3b_or3b_wx181 = multm_reduce_mulb1_add3b_maj3b_wx181 | multm_reduce_mulb1_add3b_maj3b_wy181;
  assign multm_reduce_mulb1_add3b_maj3b_wx0 = multm_reduce_mulb1_sq1 & multm_reduce_mulb1_cq0;
  assign multm_reduce_mulb1_add3b_maj3b_wx1 = multm_reduce_mulb1_sq2 & multm_reduce_mulb1_cq1;
  assign multm_reduce_mulb1_add3b_maj3b_wx4 = multm_reduce_mulb1_sq5 & multm_reduce_mulb1_cq4;
  assign multm_reduce_mulb1_add3b_maj3b_wx5 = multm_reduce_mulb1_sq6 & multm_reduce_mulb1_cq5;
  assign multm_reduce_mulb1_add3b_maj3b_wx6 = multm_reduce_mulb1_sq7 & multm_reduce_mulb1_cq6;
  assign multm_reduce_mulb1_add3b_maj3b_wx7 = multm_reduce_mulb1_sq8 & multm_reduce_mulb1_cq7;
  assign multm_reduce_mulb1_add3b_maj3b_wx10 = multm_reduce_mulb1_sq11 & multm_reduce_mulb1_cq10;
  assign multm_reduce_mulb1_add3b_maj3b_wx12 = multm_reduce_mulb1_sq13 & multm_reduce_mulb1_cq12;
  assign multm_reduce_mulb1_add3b_maj3b_wx18 = multm_reduce_mulb1_sq19 & multm_reduce_mulb1_cq18;
  assign multm_reduce_mulb1_add3b_maj3b_wx20 = multm_reduce_mulb1_sq21 & multm_reduce_mulb1_cq20;
  assign multm_reduce_mulb1_add3b_maj3b_wx22 = multm_reduce_mulb1_sq23 & multm_reduce_mulb1_cq22;
  assign multm_reduce_mulb1_add3b_maj3b_wx23 = multm_reduce_mulb1_sq24 & multm_reduce_mulb1_cq23;
  assign multm_reduce_mulb1_add3b_maj3b_wx24 = multm_reduce_mulb1_sq25 & multm_reduce_mulb1_cq24;
  assign multm_reduce_mulb1_add3b_maj3b_wx28 = multm_reduce_mulb1_sq29 & multm_reduce_mulb1_cq28;
  assign multm_reduce_mulb1_add3b_maj3b_wx30 = multm_reduce_mulb1_sq31 & multm_reduce_mulb1_cq30;
  assign multm_reduce_mulb1_add3b_maj3b_wx32 = multm_reduce_mulb1_sq33 & multm_reduce_mulb1_cq32;
  assign multm_reduce_mulb1_add3b_maj3b_wx34 = multm_reduce_mulb1_sq35 & multm_reduce_mulb1_cq34;
  assign multm_reduce_mulb1_add3b_maj3b_wx37 = multm_reduce_mulb1_sq38 & multm_reduce_mulb1_cq37;
  assign multm_reduce_mulb1_add3b_maj3b_wx40 = multm_reduce_mulb1_sq41 & multm_reduce_mulb1_cq40;
  assign multm_reduce_mulb1_add3b_maj3b_wx41 = multm_reduce_mulb1_sq42 & multm_reduce_mulb1_cq41;
  assign multm_reduce_mulb1_add3b_maj3b_wx42 = multm_reduce_mulb1_sq43 & multm_reduce_mulb1_cq42;
  assign multm_reduce_mulb1_add3b_maj3b_wx43 = multm_reduce_mulb1_sq44 & multm_reduce_mulb1_cq43;
  assign multm_reduce_mulb1_add3b_maj3b_wx47 = multm_reduce_mulb1_sq48 & multm_reduce_mulb1_cq47;
  assign multm_reduce_mulb1_add3b_maj3b_wx48 = multm_reduce_mulb1_sq49 & multm_reduce_mulb1_cq48;
  assign multm_reduce_mulb1_add3b_maj3b_wx51 = multm_reduce_mulb1_sq52 & multm_reduce_mulb1_cq51;
  assign multm_reduce_mulb1_add3b_maj3b_wx52 = multm_reduce_mulb1_sq53 & multm_reduce_mulb1_cq52;
  assign multm_reduce_mulb1_add3b_maj3b_wx53 = multm_reduce_mulb1_sq54 & multm_reduce_mulb1_cq53;
  assign multm_reduce_mulb1_add3b_maj3b_wx54 = multm_reduce_mulb1_sq55 & multm_reduce_mulb1_cq54;
  assign multm_reduce_mulb1_add3b_maj3b_wx55 = multm_reduce_mulb1_sq56 & multm_reduce_mulb1_cq55;
  assign multm_reduce_mulb1_add3b_maj3b_wx57 = multm_reduce_mulb1_sq58 & multm_reduce_mulb1_cq57;
  assign multm_reduce_mulb1_add3b_maj3b_wx62 = multm_reduce_mulb1_sq63 & multm_reduce_mulb1_cq62;
  assign multm_reduce_mulb1_add3b_maj3b_wx66 = multm_reduce_mulb1_sq67 & multm_reduce_mulb1_cq66;
  assign multm_reduce_mulb1_add3b_maj3b_wx68 = multm_reduce_mulb1_sq69 & multm_reduce_mulb1_cq68;
  assign multm_reduce_mulb1_add3b_maj3b_wx69 = multm_reduce_mulb1_sq70 & multm_reduce_mulb1_cq69;
  assign multm_reduce_mulb1_add3b_maj3b_wx71 = multm_reduce_mulb1_sq72 & multm_reduce_mulb1_cq71;
  assign multm_reduce_mulb1_add3b_maj3b_wx73 = multm_reduce_mulb1_sq74 & multm_reduce_mulb1_cq73;
  assign multm_reduce_mulb1_add3b_maj3b_wx74 = multm_reduce_mulb1_sq75 & multm_reduce_mulb1_cq74;
  assign multm_reduce_mulb1_add3b_maj3b_wx79 = multm_reduce_mulb1_sq80 & multm_reduce_mulb1_cq79;
  assign multm_reduce_mulb1_add3b_maj3b_wx80 = multm_reduce_mulb1_sq81 & multm_reduce_mulb1_cq80;
  assign multm_reduce_mulb1_add3b_maj3b_wx82 = multm_reduce_mulb1_sq83 & multm_reduce_mulb1_cq82;
  assign multm_reduce_mulb1_add3b_maj3b_wx86 = multm_reduce_mulb1_sq87 & multm_reduce_mulb1_cq86;
  assign multm_reduce_mulb1_add3b_maj3b_wx88 = multm_reduce_mulb1_sq89 & multm_reduce_mulb1_cq88;
  assign multm_reduce_mulb1_add3b_maj3b_wx90 = multm_reduce_mulb1_sq91 & multm_reduce_mulb1_cq90;
  assign multm_reduce_mulb1_add3b_maj3b_wx91 = multm_reduce_mulb1_sq92 & multm_reduce_mulb1_cq91;
  assign multm_reduce_mulb1_add3b_maj3b_wx96 = multm_reduce_mulb1_sq97 & multm_reduce_mulb1_cq96;
  assign multm_reduce_mulb1_add3b_maj3b_wx99 = multm_reduce_mulb1_sq100 & multm_reduce_mulb1_cq99;
  assign multm_reduce_mulb1_add3b_maj3b_wx100 = multm_reduce_mulb1_sq101 & multm_reduce_mulb1_cq100;
  assign multm_reduce_mulb1_add3b_maj3b_wx101 = multm_reduce_mulb1_sq102 & multm_reduce_mulb1_cq101;
  assign multm_reduce_mulb1_add3b_maj3b_wx102 = multm_reduce_mulb1_sq103 & multm_reduce_mulb1_cq102;
  assign multm_reduce_mulb1_add3b_maj3b_wx104 = multm_reduce_mulb1_sq105 & multm_reduce_mulb1_cq104;
  assign multm_reduce_mulb1_add3b_maj3b_wx105 = multm_reduce_mulb1_sq106 & multm_reduce_mulb1_cq105;
  assign multm_reduce_mulb1_add3b_maj3b_wx107 = multm_reduce_mulb1_sq108 & multm_reduce_mulb1_cq107;
  assign multm_reduce_mulb1_add3b_maj3b_wx108 = multm_reduce_mulb1_sq109 & multm_reduce_mulb1_cq108;
  assign multm_reduce_mulb1_add3b_maj3b_wx109 = multm_reduce_mulb1_sq110 & multm_reduce_mulb1_cq109;
  assign multm_reduce_mulb1_add3b_maj3b_wx110 = multm_reduce_mulb1_sq111 & multm_reduce_mulb1_cq110;
  assign multm_reduce_mulb1_add3b_maj3b_wx112 = multm_reduce_mulb1_sq113 & multm_reduce_mulb1_cq112;
  assign multm_reduce_mulb1_add3b_maj3b_wx114 = multm_reduce_mulb1_sq115 & multm_reduce_mulb1_cq114;
  assign multm_reduce_mulb1_add3b_maj3b_wx117 = multm_reduce_mulb1_sq118 & multm_reduce_mulb1_cq117;
  assign multm_reduce_mulb1_add3b_maj3b_wx118 = multm_reduce_mulb1_sq119 & multm_reduce_mulb1_cq118;
  assign multm_reduce_mulb1_add3b_maj3b_wx119 = multm_reduce_mulb1_sq120 & multm_reduce_mulb1_cq119;
  assign multm_reduce_mulb1_add3b_maj3b_wx120 = multm_reduce_mulb1_sq121 & multm_reduce_mulb1_cq120;
  assign multm_reduce_mulb1_add3b_maj3b_wx121 = multm_reduce_mulb1_sq122 & multm_reduce_mulb1_cq121;
  assign multm_reduce_mulb1_add3b_maj3b_wx122 = multm_reduce_mulb1_sq123 & multm_reduce_mulb1_cq122;
  assign multm_reduce_mulb1_add3b_maj3b_wx123 = multm_reduce_mulb1_sq124 & multm_reduce_mulb1_cq123;
  assign multm_reduce_mulb1_add3b_maj3b_wx128 = multm_reduce_mulb1_sq129 & multm_reduce_mulb1_cq128;
  assign multm_reduce_mulb1_add3b_maj3b_wx130 = multm_reduce_mulb1_sq131 & multm_reduce_mulb1_cq130;
  assign multm_reduce_mulb1_add3b_maj3b_wx132 = multm_reduce_mulb1_sq133 & multm_reduce_mulb1_cq132;
  assign multm_reduce_mulb1_add3b_maj3b_wx135 = multm_reduce_mulb1_sq136 & multm_reduce_mulb1_cq135;
  assign multm_reduce_mulb1_add3b_maj3b_wx136 = multm_reduce_mulb1_sq137 & multm_reduce_mulb1_cq136;
  assign multm_reduce_mulb1_add3b_maj3b_wx140 = multm_reduce_mulb1_sq141 & multm_reduce_mulb1_cq140;
  assign multm_reduce_mulb1_add3b_maj3b_wx141 = multm_reduce_mulb1_sq142 & multm_reduce_mulb1_cq141;
  assign multm_reduce_mulb1_add3b_maj3b_wx142 = multm_reduce_mulb1_sq143 & multm_reduce_mulb1_cq142;
  assign multm_reduce_mulb1_add3b_maj3b_wx143 = multm_reduce_mulb1_sq144 & multm_reduce_mulb1_cq143;
  assign multm_reduce_mulb1_add3b_maj3b_wx144 = multm_reduce_mulb1_sq145 & multm_reduce_mulb1_cq144;
  assign multm_reduce_mulb1_add3b_maj3b_wx147 = multm_reduce_mulb1_sq148 & multm_reduce_mulb1_cq147;
  assign multm_reduce_mulb1_add3b_maj3b_wx150 = multm_reduce_mulb1_sq151 & multm_reduce_mulb1_cq150;
  assign multm_reduce_mulb1_add3b_maj3b_wx151 = multm_reduce_mulb1_sq152 & multm_reduce_mulb1_cq151;
  assign multm_reduce_mulb1_add3b_maj3b_wx152 = multm_reduce_mulb1_sq153 & multm_reduce_mulb1_cq152;
  assign multm_reduce_mulb1_add3b_maj3b_wx153 = multm_reduce_mulb1_sq154 & multm_reduce_mulb1_cq153;
  assign multm_reduce_mulb1_add3b_maj3b_wx155 = multm_reduce_mulb1_sq156 & multm_reduce_mulb1_cq155;
  assign multm_reduce_mulb1_add3b_maj3b_wx156 = multm_reduce_mulb1_sq157 & multm_reduce_mulb1_cq156;
  assign multm_reduce_mulb1_add3b_maj3b_wx157 = multm_reduce_mulb1_sq158 & multm_reduce_mulb1_cq157;
  assign multm_reduce_mulb1_add3b_maj3b_wx158 = multm_reduce_mulb1_sq159 & multm_reduce_mulb1_cq158;
  assign multm_reduce_mulb1_add3b_maj3b_wx159 = multm_reduce_mulb1_sq160 & multm_reduce_mulb1_cq159;
  assign multm_reduce_mulb1_add3b_maj3b_wx160 = multm_reduce_mulb1_sq161 & multm_reduce_mulb1_cq160;
  assign multm_reduce_mulb1_add3b_maj3b_wx162 = multm_reduce_mulb1_sq163 & multm_reduce_mulb1_cq162;
  assign multm_reduce_mulb1_add3b_maj3b_wx166 = multm_reduce_mulb1_sq167 & multm_reduce_mulb1_cq166;
  assign multm_reduce_mulb1_add3b_maj3b_wx171 = multm_reduce_mulb1_sq172 & multm_reduce_mulb1_cq171;
  assign multm_reduce_mulb1_add3b_maj3b_wx172 = multm_reduce_mulb1_sq173 & multm_reduce_mulb1_cq172;
  assign multm_reduce_mulb1_add3b_maj3b_wx173 = multm_reduce_mulb1_sq174 & multm_reduce_mulb1_cq173;
  assign multm_reduce_mulb1_add3b_maj3b_wx174 = multm_reduce_mulb1_sq175 & multm_reduce_mulb1_cq174;
  assign multm_reduce_mulb1_add3b_maj3b_wx175 = multm_reduce_mulb1_sq176 & multm_reduce_mulb1_cq175;
  assign multm_reduce_mulb1_add3b_maj3b_wx179 = multm_reduce_mulb1_sq180 & multm_reduce_mulb1_cq179;
  assign multm_reduce_mulb1_add3b_maj3b_wx181 = multm_reduce_mulb1_sq182 & multm_reduce_mulb1_cq181;
  assign multm_reduce_mulb1_add3b_maj3b_wy0 = multm_reduce_mulb1_sq1 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy1 = multm_reduce_mulb1_sq2 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy4 = multm_reduce_mulb1_sq5 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy5 = multm_reduce_mulb1_sq6 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy6 = multm_reduce_mulb1_sq7 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy7 = multm_reduce_mulb1_sq8 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy10 = multm_reduce_mulb1_sq11 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy12 = multm_reduce_mulb1_sq13 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy18 = multm_reduce_mulb1_sq19 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy20 = multm_reduce_mulb1_sq21 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy22 = multm_reduce_mulb1_sq23 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy23 = multm_reduce_mulb1_sq24 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy24 = multm_reduce_mulb1_sq25 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy28 = multm_reduce_mulb1_sq29 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy30 = multm_reduce_mulb1_sq31 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy32 = multm_reduce_mulb1_sq33 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy34 = multm_reduce_mulb1_sq35 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy37 = multm_reduce_mulb1_sq38 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy40 = multm_reduce_mulb1_sq41 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy41 = multm_reduce_mulb1_sq42 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy42 = multm_reduce_mulb1_sq43 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy43 = multm_reduce_mulb1_sq44 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy47 = multm_reduce_mulb1_sq48 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy48 = multm_reduce_mulb1_sq49 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy51 = multm_reduce_mulb1_sq52 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy52 = multm_reduce_mulb1_sq53 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy53 = multm_reduce_mulb1_sq54 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy54 = multm_reduce_mulb1_sq55 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy55 = multm_reduce_mulb1_sq56 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy57 = multm_reduce_mulb1_sq58 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy62 = multm_reduce_mulb1_sq63 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy66 = multm_reduce_mulb1_sq67 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy68 = multm_reduce_mulb1_sq69 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy69 = multm_reduce_mulb1_sq70 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy71 = multm_reduce_mulb1_sq72 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy73 = multm_reduce_mulb1_sq74 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy74 = multm_reduce_mulb1_sq75 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy79 = multm_reduce_mulb1_sq80 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy80 = multm_reduce_mulb1_sq81 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy82 = multm_reduce_mulb1_sq83 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy86 = multm_reduce_mulb1_sq87 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy88 = multm_reduce_mulb1_sq89 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy90 = multm_reduce_mulb1_sq91 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy91 = multm_reduce_mulb1_sq92 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy96 = multm_reduce_mulb1_sq97 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy99 = multm_reduce_mulb1_sq100 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy100 = multm_reduce_mulb1_sq101 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy101 = multm_reduce_mulb1_sq102 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy102 = multm_reduce_mulb1_sq103 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy104 = multm_reduce_mulb1_sq105 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy105 = multm_reduce_mulb1_sq106 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy107 = multm_reduce_mulb1_sq108 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy108 = multm_reduce_mulb1_sq109 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy109 = multm_reduce_mulb1_sq110 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy110 = multm_reduce_mulb1_sq111 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy112 = multm_reduce_mulb1_sq113 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy114 = multm_reduce_mulb1_sq115 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy117 = multm_reduce_mulb1_sq118 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy118 = multm_reduce_mulb1_sq119 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy119 = multm_reduce_mulb1_sq120 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy120 = multm_reduce_mulb1_sq121 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy121 = multm_reduce_mulb1_sq122 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy122 = multm_reduce_mulb1_sq123 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy123 = multm_reduce_mulb1_sq124 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy128 = multm_reduce_mulb1_sq129 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy130 = multm_reduce_mulb1_sq131 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy132 = multm_reduce_mulb1_sq133 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy135 = multm_reduce_mulb1_sq136 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy136 = multm_reduce_mulb1_sq137 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy140 = multm_reduce_mulb1_sq141 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy141 = multm_reduce_mulb1_sq142 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy142 = multm_reduce_mulb1_sq143 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy143 = multm_reduce_mulb1_sq144 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy144 = multm_reduce_mulb1_sq145 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy147 = multm_reduce_mulb1_sq148 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy150 = multm_reduce_mulb1_sq151 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy151 = multm_reduce_mulb1_sq152 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy152 = multm_reduce_mulb1_sq153 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy153 = multm_reduce_mulb1_sq154 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy155 = multm_reduce_mulb1_sq156 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy156 = multm_reduce_mulb1_sq157 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy157 = multm_reduce_mulb1_sq158 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy158 = multm_reduce_mulb1_sq159 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy159 = multm_reduce_mulb1_sq160 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy160 = multm_reduce_mulb1_sq161 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy162 = multm_reduce_mulb1_sq163 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy166 = multm_reduce_mulb1_sq167 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy171 = multm_reduce_mulb1_sq172 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy172 = multm_reduce_mulb1_sq173 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy173 = multm_reduce_mulb1_sq174 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy174 = multm_reduce_mulb1_sq175 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy175 = multm_reduce_mulb1_sq176 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy179 = multm_reduce_mulb1_sq180 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_wy181 = multm_reduce_mulb1_sq182 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy0 = multm_reduce_mulb1_cq0 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy1 = multm_reduce_mulb1_cq1 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy4 = multm_reduce_mulb1_cq4 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy5 = multm_reduce_mulb1_cq5 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy6 = multm_reduce_mulb1_cq6 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy7 = multm_reduce_mulb1_cq7 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy10 = multm_reduce_mulb1_cq10 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy12 = multm_reduce_mulb1_cq12 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy18 = multm_reduce_mulb1_cq18 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy20 = multm_reduce_mulb1_cq20 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy22 = multm_reduce_mulb1_cq22 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy23 = multm_reduce_mulb1_cq23 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy24 = multm_reduce_mulb1_cq24 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy28 = multm_reduce_mulb1_cq28 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy30 = multm_reduce_mulb1_cq30 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy32 = multm_reduce_mulb1_cq32 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy34 = multm_reduce_mulb1_cq34 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy37 = multm_reduce_mulb1_cq37 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy40 = multm_reduce_mulb1_cq40 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy41 = multm_reduce_mulb1_cq41 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy42 = multm_reduce_mulb1_cq42 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy43 = multm_reduce_mulb1_cq43 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy47 = multm_reduce_mulb1_cq47 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy48 = multm_reduce_mulb1_cq48 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy51 = multm_reduce_mulb1_cq51 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy52 = multm_reduce_mulb1_cq52 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy53 = multm_reduce_mulb1_cq53 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy54 = multm_reduce_mulb1_cq54 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy55 = multm_reduce_mulb1_cq55 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy57 = multm_reduce_mulb1_cq57 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy62 = multm_reduce_mulb1_cq62 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy66 = multm_reduce_mulb1_cq66 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy68 = multm_reduce_mulb1_cq68 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy69 = multm_reduce_mulb1_cq69 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy71 = multm_reduce_mulb1_cq71 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy73 = multm_reduce_mulb1_cq73 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy74 = multm_reduce_mulb1_cq74 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy79 = multm_reduce_mulb1_cq79 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy80 = multm_reduce_mulb1_cq80 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy82 = multm_reduce_mulb1_cq82 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy86 = multm_reduce_mulb1_cq86 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy88 = multm_reduce_mulb1_cq88 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy90 = multm_reduce_mulb1_cq90 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy91 = multm_reduce_mulb1_cq91 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy96 = multm_reduce_mulb1_cq96 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy99 = multm_reduce_mulb1_cq99 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy100 = multm_reduce_mulb1_cq100 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy101 = multm_reduce_mulb1_cq101 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy102 = multm_reduce_mulb1_cq102 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy104 = multm_reduce_mulb1_cq104 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy105 = multm_reduce_mulb1_cq105 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy107 = multm_reduce_mulb1_cq107 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy108 = multm_reduce_mulb1_cq108 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy109 = multm_reduce_mulb1_cq109 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy110 = multm_reduce_mulb1_cq110 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy112 = multm_reduce_mulb1_cq112 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy114 = multm_reduce_mulb1_cq114 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy117 = multm_reduce_mulb1_cq117 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy118 = multm_reduce_mulb1_cq118 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy119 = multm_reduce_mulb1_cq119 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy120 = multm_reduce_mulb1_cq120 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy121 = multm_reduce_mulb1_cq121 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy122 = multm_reduce_mulb1_cq122 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy123 = multm_reduce_mulb1_cq123 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy128 = multm_reduce_mulb1_cq128 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy130 = multm_reduce_mulb1_cq130 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy132 = multm_reduce_mulb1_cq132 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy135 = multm_reduce_mulb1_cq135 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy136 = multm_reduce_mulb1_cq136 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy140 = multm_reduce_mulb1_cq140 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy141 = multm_reduce_mulb1_cq141 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy142 = multm_reduce_mulb1_cq142 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy143 = multm_reduce_mulb1_cq143 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy144 = multm_reduce_mulb1_cq144 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy147 = multm_reduce_mulb1_cq147 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy150 = multm_reduce_mulb1_cq150 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy151 = multm_reduce_mulb1_cq151 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy152 = multm_reduce_mulb1_cq152 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy153 = multm_reduce_mulb1_cq153 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy155 = multm_reduce_mulb1_cq155 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy156 = multm_reduce_mulb1_cq156 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy157 = multm_reduce_mulb1_cq157 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy158 = multm_reduce_mulb1_cq158 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy159 = multm_reduce_mulb1_cq159 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy160 = multm_reduce_mulb1_cq160 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy162 = multm_reduce_mulb1_cq162 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy166 = multm_reduce_mulb1_cq166 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy171 = multm_reduce_mulb1_cq171 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy172 = multm_reduce_mulb1_cq172 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy173 = multm_reduce_mulb1_cq173 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy174 = multm_reduce_mulb1_cq174 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy175 = multm_reduce_mulb1_cq175 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy179 = multm_reduce_mulb1_cq179 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_maj3b_xy181 = multm_reduce_mulb1_cq181 & multm_reduce_qb2;
  assign multm_reduce_mulb1_add3b_xor3b_wx0 = multm_reduce_mulb1_sq1 ^ multm_reduce_mulb1_cq0;
  assign multm_reduce_mulb1_add3b_xor3b_wx1 = multm_reduce_mulb1_sq2 ^ multm_reduce_mulb1_cq1;
  assign multm_reduce_mulb1_add3b_xor3b_wx4 = multm_reduce_mulb1_sq5 ^ multm_reduce_mulb1_cq4;
  assign multm_reduce_mulb1_add3b_xor3b_wx5 = multm_reduce_mulb1_sq6 ^ multm_reduce_mulb1_cq5;
  assign multm_reduce_mulb1_add3b_xor3b_wx6 = multm_reduce_mulb1_sq7 ^ multm_reduce_mulb1_cq6;
  assign multm_reduce_mulb1_add3b_xor3b_wx7 = multm_reduce_mulb1_sq8 ^ multm_reduce_mulb1_cq7;
  assign multm_reduce_mulb1_add3b_xor3b_wx10 = multm_reduce_mulb1_sq11 ^ multm_reduce_mulb1_cq10;
  assign multm_reduce_mulb1_add3b_xor3b_wx12 = multm_reduce_mulb1_sq13 ^ multm_reduce_mulb1_cq12;
  assign multm_reduce_mulb1_add3b_xor3b_wx18 = multm_reduce_mulb1_sq19 ^ multm_reduce_mulb1_cq18;
  assign multm_reduce_mulb1_add3b_xor3b_wx20 = multm_reduce_mulb1_sq21 ^ multm_reduce_mulb1_cq20;
  assign multm_reduce_mulb1_add3b_xor3b_wx22 = multm_reduce_mulb1_sq23 ^ multm_reduce_mulb1_cq22;
  assign multm_reduce_mulb1_add3b_xor3b_wx23 = multm_reduce_mulb1_sq24 ^ multm_reduce_mulb1_cq23;
  assign multm_reduce_mulb1_add3b_xor3b_wx24 = multm_reduce_mulb1_sq25 ^ multm_reduce_mulb1_cq24;
  assign multm_reduce_mulb1_add3b_xor3b_wx28 = multm_reduce_mulb1_sq29 ^ multm_reduce_mulb1_cq28;
  assign multm_reduce_mulb1_add3b_xor3b_wx30 = multm_reduce_mulb1_sq31 ^ multm_reduce_mulb1_cq30;
  assign multm_reduce_mulb1_add3b_xor3b_wx32 = multm_reduce_mulb1_sq33 ^ multm_reduce_mulb1_cq32;
  assign multm_reduce_mulb1_add3b_xor3b_wx34 = multm_reduce_mulb1_sq35 ^ multm_reduce_mulb1_cq34;
  assign multm_reduce_mulb1_add3b_xor3b_wx37 = multm_reduce_mulb1_sq38 ^ multm_reduce_mulb1_cq37;
  assign multm_reduce_mulb1_add3b_xor3b_wx40 = multm_reduce_mulb1_sq41 ^ multm_reduce_mulb1_cq40;
  assign multm_reduce_mulb1_add3b_xor3b_wx41 = multm_reduce_mulb1_sq42 ^ multm_reduce_mulb1_cq41;
  assign multm_reduce_mulb1_add3b_xor3b_wx42 = multm_reduce_mulb1_sq43 ^ multm_reduce_mulb1_cq42;
  assign multm_reduce_mulb1_add3b_xor3b_wx43 = multm_reduce_mulb1_sq44 ^ multm_reduce_mulb1_cq43;
  assign multm_reduce_mulb1_add3b_xor3b_wx47 = multm_reduce_mulb1_sq48 ^ multm_reduce_mulb1_cq47;
  assign multm_reduce_mulb1_add3b_xor3b_wx48 = multm_reduce_mulb1_sq49 ^ multm_reduce_mulb1_cq48;
  assign multm_reduce_mulb1_add3b_xor3b_wx51 = multm_reduce_mulb1_sq52 ^ multm_reduce_mulb1_cq51;
  assign multm_reduce_mulb1_add3b_xor3b_wx52 = multm_reduce_mulb1_sq53 ^ multm_reduce_mulb1_cq52;
  assign multm_reduce_mulb1_add3b_xor3b_wx53 = multm_reduce_mulb1_sq54 ^ multm_reduce_mulb1_cq53;
  assign multm_reduce_mulb1_add3b_xor3b_wx54 = multm_reduce_mulb1_sq55 ^ multm_reduce_mulb1_cq54;
  assign multm_reduce_mulb1_add3b_xor3b_wx55 = multm_reduce_mulb1_sq56 ^ multm_reduce_mulb1_cq55;
  assign multm_reduce_mulb1_add3b_xor3b_wx57 = multm_reduce_mulb1_sq58 ^ multm_reduce_mulb1_cq57;
  assign multm_reduce_mulb1_add3b_xor3b_wx62 = multm_reduce_mulb1_sq63 ^ multm_reduce_mulb1_cq62;
  assign multm_reduce_mulb1_add3b_xor3b_wx66 = multm_reduce_mulb1_sq67 ^ multm_reduce_mulb1_cq66;
  assign multm_reduce_mulb1_add3b_xor3b_wx68 = multm_reduce_mulb1_sq69 ^ multm_reduce_mulb1_cq68;
  assign multm_reduce_mulb1_add3b_xor3b_wx69 = multm_reduce_mulb1_sq70 ^ multm_reduce_mulb1_cq69;
  assign multm_reduce_mulb1_add3b_xor3b_wx71 = multm_reduce_mulb1_sq72 ^ multm_reduce_mulb1_cq71;
  assign multm_reduce_mulb1_add3b_xor3b_wx73 = multm_reduce_mulb1_sq74 ^ multm_reduce_mulb1_cq73;
  assign multm_reduce_mulb1_add3b_xor3b_wx74 = multm_reduce_mulb1_sq75 ^ multm_reduce_mulb1_cq74;
  assign multm_reduce_mulb1_add3b_xor3b_wx79 = multm_reduce_mulb1_sq80 ^ multm_reduce_mulb1_cq79;
  assign multm_reduce_mulb1_add3b_xor3b_wx80 = multm_reduce_mulb1_sq81 ^ multm_reduce_mulb1_cq80;
  assign multm_reduce_mulb1_add3b_xor3b_wx82 = multm_reduce_mulb1_sq83 ^ multm_reduce_mulb1_cq82;
  assign multm_reduce_mulb1_add3b_xor3b_wx86 = multm_reduce_mulb1_sq87 ^ multm_reduce_mulb1_cq86;
  assign multm_reduce_mulb1_add3b_xor3b_wx88 = multm_reduce_mulb1_sq89 ^ multm_reduce_mulb1_cq88;
  assign multm_reduce_mulb1_add3b_xor3b_wx90 = multm_reduce_mulb1_sq91 ^ multm_reduce_mulb1_cq90;
  assign multm_reduce_mulb1_add3b_xor3b_wx91 = multm_reduce_mulb1_sq92 ^ multm_reduce_mulb1_cq91;
  assign multm_reduce_mulb1_add3b_xor3b_wx96 = multm_reduce_mulb1_sq97 ^ multm_reduce_mulb1_cq96;
  assign multm_reduce_mulb1_add3b_xor3b_wx99 = multm_reduce_mulb1_sq100 ^ multm_reduce_mulb1_cq99;
  assign multm_reduce_mulb1_add3b_xor3b_wx100 = multm_reduce_mulb1_sq101 ^ multm_reduce_mulb1_cq100;
  assign multm_reduce_mulb1_add3b_xor3b_wx101 = multm_reduce_mulb1_sq102 ^ multm_reduce_mulb1_cq101;
  assign multm_reduce_mulb1_add3b_xor3b_wx102 = multm_reduce_mulb1_sq103 ^ multm_reduce_mulb1_cq102;
  assign multm_reduce_mulb1_add3b_xor3b_wx104 = multm_reduce_mulb1_sq105 ^ multm_reduce_mulb1_cq104;
  assign multm_reduce_mulb1_add3b_xor3b_wx105 = multm_reduce_mulb1_sq106 ^ multm_reduce_mulb1_cq105;
  assign multm_reduce_mulb1_add3b_xor3b_wx107 = multm_reduce_mulb1_sq108 ^ multm_reduce_mulb1_cq107;
  assign multm_reduce_mulb1_add3b_xor3b_wx108 = multm_reduce_mulb1_sq109 ^ multm_reduce_mulb1_cq108;
  assign multm_reduce_mulb1_add3b_xor3b_wx109 = multm_reduce_mulb1_sq110 ^ multm_reduce_mulb1_cq109;
  assign multm_reduce_mulb1_add3b_xor3b_wx110 = multm_reduce_mulb1_sq111 ^ multm_reduce_mulb1_cq110;
  assign multm_reduce_mulb1_add3b_xor3b_wx112 = multm_reduce_mulb1_sq113 ^ multm_reduce_mulb1_cq112;
  assign multm_reduce_mulb1_add3b_xor3b_wx114 = multm_reduce_mulb1_sq115 ^ multm_reduce_mulb1_cq114;
  assign multm_reduce_mulb1_add3b_xor3b_wx117 = multm_reduce_mulb1_sq118 ^ multm_reduce_mulb1_cq117;
  assign multm_reduce_mulb1_add3b_xor3b_wx118 = multm_reduce_mulb1_sq119 ^ multm_reduce_mulb1_cq118;
  assign multm_reduce_mulb1_add3b_xor3b_wx119 = multm_reduce_mulb1_sq120 ^ multm_reduce_mulb1_cq119;
  assign multm_reduce_mulb1_add3b_xor3b_wx120 = multm_reduce_mulb1_sq121 ^ multm_reduce_mulb1_cq120;
  assign multm_reduce_mulb1_add3b_xor3b_wx121 = multm_reduce_mulb1_sq122 ^ multm_reduce_mulb1_cq121;
  assign multm_reduce_mulb1_add3b_xor3b_wx122 = multm_reduce_mulb1_sq123 ^ multm_reduce_mulb1_cq122;
  assign multm_reduce_mulb1_add3b_xor3b_wx123 = multm_reduce_mulb1_sq124 ^ multm_reduce_mulb1_cq123;
  assign multm_reduce_mulb1_add3b_xor3b_wx128 = multm_reduce_mulb1_sq129 ^ multm_reduce_mulb1_cq128;
  assign multm_reduce_mulb1_add3b_xor3b_wx130 = multm_reduce_mulb1_sq131 ^ multm_reduce_mulb1_cq130;
  assign multm_reduce_mulb1_add3b_xor3b_wx132 = multm_reduce_mulb1_sq133 ^ multm_reduce_mulb1_cq132;
  assign multm_reduce_mulb1_add3b_xor3b_wx135 = multm_reduce_mulb1_sq136 ^ multm_reduce_mulb1_cq135;
  assign multm_reduce_mulb1_add3b_xor3b_wx136 = multm_reduce_mulb1_sq137 ^ multm_reduce_mulb1_cq136;
  assign multm_reduce_mulb1_add3b_xor3b_wx140 = multm_reduce_mulb1_sq141 ^ multm_reduce_mulb1_cq140;
  assign multm_reduce_mulb1_add3b_xor3b_wx141 = multm_reduce_mulb1_sq142 ^ multm_reduce_mulb1_cq141;
  assign multm_reduce_mulb1_add3b_xor3b_wx142 = multm_reduce_mulb1_sq143 ^ multm_reduce_mulb1_cq142;
  assign multm_reduce_mulb1_add3b_xor3b_wx143 = multm_reduce_mulb1_sq144 ^ multm_reduce_mulb1_cq143;
  assign multm_reduce_mulb1_add3b_xor3b_wx144 = multm_reduce_mulb1_sq145 ^ multm_reduce_mulb1_cq144;
  assign multm_reduce_mulb1_add3b_xor3b_wx147 = multm_reduce_mulb1_sq148 ^ multm_reduce_mulb1_cq147;
  assign multm_reduce_mulb1_add3b_xor3b_wx150 = multm_reduce_mulb1_sq151 ^ multm_reduce_mulb1_cq150;
  assign multm_reduce_mulb1_add3b_xor3b_wx151 = multm_reduce_mulb1_sq152 ^ multm_reduce_mulb1_cq151;
  assign multm_reduce_mulb1_add3b_xor3b_wx152 = multm_reduce_mulb1_sq153 ^ multm_reduce_mulb1_cq152;
  assign multm_reduce_mulb1_add3b_xor3b_wx153 = multm_reduce_mulb1_sq154 ^ multm_reduce_mulb1_cq153;
  assign multm_reduce_mulb1_add3b_xor3b_wx155 = multm_reduce_mulb1_sq156 ^ multm_reduce_mulb1_cq155;
  assign multm_reduce_mulb1_add3b_xor3b_wx156 = multm_reduce_mulb1_sq157 ^ multm_reduce_mulb1_cq156;
  assign multm_reduce_mulb1_add3b_xor3b_wx157 = multm_reduce_mulb1_sq158 ^ multm_reduce_mulb1_cq157;
  assign multm_reduce_mulb1_add3b_xor3b_wx158 = multm_reduce_mulb1_sq159 ^ multm_reduce_mulb1_cq158;
  assign multm_reduce_mulb1_add3b_xor3b_wx159 = multm_reduce_mulb1_sq160 ^ multm_reduce_mulb1_cq159;
  assign multm_reduce_mulb1_add3b_xor3b_wx160 = multm_reduce_mulb1_sq161 ^ multm_reduce_mulb1_cq160;
  assign multm_reduce_mulb1_add3b_xor3b_wx162 = multm_reduce_mulb1_sq163 ^ multm_reduce_mulb1_cq162;
  assign multm_reduce_mulb1_add3b_xor3b_wx166 = multm_reduce_mulb1_sq167 ^ multm_reduce_mulb1_cq166;
  assign multm_reduce_mulb1_add3b_xor3b_wx171 = multm_reduce_mulb1_sq172 ^ multm_reduce_mulb1_cq171;
  assign multm_reduce_mulb1_add3b_xor3b_wx172 = multm_reduce_mulb1_sq173 ^ multm_reduce_mulb1_cq172;
  assign multm_reduce_mulb1_add3b_xor3b_wx173 = multm_reduce_mulb1_sq174 ^ multm_reduce_mulb1_cq173;
  assign multm_reduce_mulb1_add3b_xor3b_wx174 = multm_reduce_mulb1_sq175 ^ multm_reduce_mulb1_cq174;
  assign multm_reduce_mulb1_add3b_xor3b_wx175 = multm_reduce_mulb1_sq176 ^ multm_reduce_mulb1_cq175;
  assign multm_reduce_mulb1_add3b_xor3b_wx179 = multm_reduce_mulb1_sq180 ^ multm_reduce_mulb1_cq179;
  assign multm_reduce_mulb1_add3b_xor3b_wx181 = multm_reduce_mulb1_sq182 ^ multm_reduce_mulb1_cq181;
  assign multm_reduce_mulb1_cq0 = xn2 & multm_reduce_sd1;
  assign multm_reduce_mulb1_cq1 = xn2 & multm_reduce_sd2;
  assign multm_reduce_mulb1_cq2 = xn2 & multm_reduce_sd3;
  assign multm_reduce_mulb1_cq3 = xn2 & multm_reduce_sd4;
  assign multm_reduce_mulb1_cq4 = xn2 & multm_reduce_sd5;
  assign multm_reduce_mulb1_cq5 = xn2 & multm_reduce_sd6;
  assign multm_reduce_mulb1_cq6 = xn2 & multm_reduce_sd7;
  assign multm_reduce_mulb1_cq7 = xn2 & multm_reduce_sd8;
  assign multm_reduce_mulb1_cq8 = xn2 & multm_reduce_sd9;
  assign multm_reduce_mulb1_cq9 = xn2 & multm_reduce_sd10;
  assign multm_reduce_mulb1_cq10 = xn2 & multm_reduce_sd11;
  assign multm_reduce_mulb1_cq11 = xn2 & multm_reduce_sd12;
  assign multm_reduce_mulb1_cq12 = xn2 & multm_reduce_sd13;
  assign multm_reduce_mulb1_cq13 = xn2 & multm_reduce_sd14;
  assign multm_reduce_mulb1_cq14 = xn2 & multm_reduce_sd15;
  assign multm_reduce_mulb1_cq15 = xn2 & multm_reduce_sd16;
  assign multm_reduce_mulb1_cq16 = xn2 & multm_reduce_sd17;
  assign multm_reduce_mulb1_cq17 = xn2 & multm_reduce_sd18;
  assign multm_reduce_mulb1_cq18 = xn2 & multm_reduce_sd19;
  assign multm_reduce_mulb1_cq19 = xn2 & multm_reduce_sd20;
  assign multm_reduce_mulb1_cq20 = xn2 & multm_reduce_sd21;
  assign multm_reduce_mulb1_cq21 = xn2 & multm_reduce_sd22;
  assign multm_reduce_mulb1_cq22 = xn2 & multm_reduce_sd23;
  assign multm_reduce_mulb1_cq23 = xn2 & multm_reduce_sd24;
  assign multm_reduce_mulb1_cq24 = xn2 & multm_reduce_sd25;
  assign multm_reduce_mulb1_cq25 = xn2 & multm_reduce_sd26;
  assign multm_reduce_mulb1_cq26 = xn2 & multm_reduce_sd27;
  assign multm_reduce_mulb1_cq27 = xn2 & multm_reduce_sd28;
  assign multm_reduce_mulb1_cq28 = xn2 & multm_reduce_sd29;
  assign multm_reduce_mulb1_cq29 = xn2 & multm_reduce_sd30;
  assign multm_reduce_mulb1_cq30 = xn2 & multm_reduce_sd31;
  assign multm_reduce_mulb1_cq31 = xn2 & multm_reduce_sd32;
  assign multm_reduce_mulb1_cq32 = xn2 & multm_reduce_sd33;
  assign multm_reduce_mulb1_cq33 = xn2 & multm_reduce_sd34;
  assign multm_reduce_mulb1_cq34 = xn2 & multm_reduce_sd35;
  assign multm_reduce_mulb1_cq35 = xn2 & multm_reduce_sd36;
  assign multm_reduce_mulb1_cq36 = xn2 & multm_reduce_sd37;
  assign multm_reduce_mulb1_cq37 = xn2 & multm_reduce_sd38;
  assign multm_reduce_mulb1_cq38 = xn2 & multm_reduce_sd39;
  assign multm_reduce_mulb1_cq39 = xn2 & multm_reduce_sd40;
  assign multm_reduce_mulb1_cq40 = xn2 & multm_reduce_sd41;
  assign multm_reduce_mulb1_cq41 = xn2 & multm_reduce_sd42;
  assign multm_reduce_mulb1_cq42 = xn2 & multm_reduce_sd43;
  assign multm_reduce_mulb1_cq43 = xn2 & multm_reduce_sd44;
  assign multm_reduce_mulb1_cq44 = xn2 & multm_reduce_sd45;
  assign multm_reduce_mulb1_cq45 = xn2 & multm_reduce_sd46;
  assign multm_reduce_mulb1_cq46 = xn2 & multm_reduce_sd47;
  assign multm_reduce_mulb1_cq47 = xn2 & multm_reduce_sd48;
  assign multm_reduce_mulb1_cq48 = xn2 & multm_reduce_sd49;
  assign multm_reduce_mulb1_cq49 = xn2 & multm_reduce_sd50;
  assign multm_reduce_mulb1_cq50 = xn2 & multm_reduce_sd51;
  assign multm_reduce_mulb1_cq51 = xn2 & multm_reduce_sd52;
  assign multm_reduce_mulb1_cq52 = xn2 & multm_reduce_sd53;
  assign multm_reduce_mulb1_cq53 = xn2 & multm_reduce_sd54;
  assign multm_reduce_mulb1_cq54 = xn2 & multm_reduce_sd55;
  assign multm_reduce_mulb1_cq55 = xn2 & multm_reduce_sd56;
  assign multm_reduce_mulb1_cq56 = xn2 & multm_reduce_sd57;
  assign multm_reduce_mulb1_cq57 = xn2 & multm_reduce_sd58;
  assign multm_reduce_mulb1_cq58 = xn2 & multm_reduce_sd59;
  assign multm_reduce_mulb1_cq59 = xn2 & multm_reduce_sd60;
  assign multm_reduce_mulb1_cq60 = xn2 & multm_reduce_sd61;
  assign multm_reduce_mulb1_cq61 = xn2 & multm_reduce_sd62;
  assign multm_reduce_mulb1_cq62 = xn2 & multm_reduce_sd63;
  assign multm_reduce_mulb1_cq63 = xn2 & multm_reduce_sd64;
  assign multm_reduce_mulb1_cq64 = xn2 & multm_reduce_sd65;
  assign multm_reduce_mulb1_cq65 = xn2 & multm_reduce_sd66;
  assign multm_reduce_mulb1_cq66 = xn2 & multm_reduce_sd67;
  assign multm_reduce_mulb1_cq67 = xn2 & multm_reduce_sd68;
  assign multm_reduce_mulb1_cq68 = xn2 & multm_reduce_sd69;
  assign multm_reduce_mulb1_cq69 = xn2 & multm_reduce_sd70;
  assign multm_reduce_mulb1_cq70 = xn2 & multm_reduce_sd71;
  assign multm_reduce_mulb1_cq71 = xn2 & multm_reduce_sd72;
  assign multm_reduce_mulb1_cq72 = xn2 & multm_reduce_sd73;
  assign multm_reduce_mulb1_cq73 = xn2 & multm_reduce_sd74;
  assign multm_reduce_mulb1_cq74 = xn2 & multm_reduce_sd75;
  assign multm_reduce_mulb1_cq75 = xn2 & multm_reduce_sd76;
  assign multm_reduce_mulb1_cq76 = xn2 & multm_reduce_sd77;
  assign multm_reduce_mulb1_cq77 = xn2 & multm_reduce_sd78;
  assign multm_reduce_mulb1_cq78 = xn2 & multm_reduce_sd79;
  assign multm_reduce_mulb1_cq79 = xn2 & multm_reduce_sd80;
  assign multm_reduce_mulb1_cq80 = xn2 & multm_reduce_sd81;
  assign multm_reduce_mulb1_cq81 = xn2 & multm_reduce_sd82;
  assign multm_reduce_mulb1_cq82 = xn2 & multm_reduce_sd83;
  assign multm_reduce_mulb1_cq83 = xn2 & multm_reduce_sd84;
  assign multm_reduce_mulb1_cq84 = xn2 & multm_reduce_sd85;
  assign multm_reduce_mulb1_cq85 = xn2 & multm_reduce_sd86;
  assign multm_reduce_mulb1_cq86 = xn2 & multm_reduce_sd87;
  assign multm_reduce_mulb1_cq87 = xn2 & multm_reduce_sd88;
  assign multm_reduce_mulb1_cq88 = xn2 & multm_reduce_sd89;
  assign multm_reduce_mulb1_cq89 = xn2 & multm_reduce_sd90;
  assign multm_reduce_mulb1_cq90 = xn2 & multm_reduce_sd91;
  assign multm_reduce_mulb1_cq91 = xn2 & multm_reduce_sd92;
  assign multm_reduce_mulb1_cq92 = xn2 & multm_reduce_sd93;
  assign multm_reduce_mulb1_cq93 = xn2 & multm_reduce_sd94;
  assign multm_reduce_mulb1_cq94 = xn2 & multm_reduce_sd95;
  assign multm_reduce_mulb1_cq95 = xn2 & multm_reduce_sd96;
  assign multm_reduce_mulb1_cq96 = xn2 & multm_reduce_sd97;
  assign multm_reduce_mulb1_cq97 = xn2 & multm_reduce_sd98;
  assign multm_reduce_mulb1_cq98 = xn2 & multm_reduce_sd99;
  assign multm_reduce_mulb1_cq99 = xn2 & multm_reduce_sd100;
  assign multm_reduce_mulb1_cq100 = xn2 & multm_reduce_sd101;
  assign multm_reduce_mulb1_cq101 = xn2 & multm_reduce_sd102;
  assign multm_reduce_mulb1_cq102 = xn2 & multm_reduce_sd103;
  assign multm_reduce_mulb1_cq103 = xn2 & multm_reduce_sd104;
  assign multm_reduce_mulb1_cq104 = xn2 & multm_reduce_sd105;
  assign multm_reduce_mulb1_cq105 = xn2 & multm_reduce_sd106;
  assign multm_reduce_mulb1_cq106 = xn2 & multm_reduce_sd107;
  assign multm_reduce_mulb1_cq107 = xn2 & multm_reduce_sd108;
  assign multm_reduce_mulb1_cq108 = xn2 & multm_reduce_sd109;
  assign multm_reduce_mulb1_cq109 = xn2 & multm_reduce_sd110;
  assign multm_reduce_mulb1_cq110 = xn2 & multm_reduce_sd111;
  assign multm_reduce_mulb1_cq111 = xn2 & multm_reduce_sd112;
  assign multm_reduce_mulb1_cq112 = xn2 & multm_reduce_sd113;
  assign multm_reduce_mulb1_cq113 = xn2 & multm_reduce_sd114;
  assign multm_reduce_mulb1_cq114 = xn2 & multm_reduce_sd115;
  assign multm_reduce_mulb1_cq115 = xn2 & multm_reduce_sd116;
  assign multm_reduce_mulb1_cq116 = xn2 & multm_reduce_sd117;
  assign multm_reduce_mulb1_cq117 = xn2 & multm_reduce_sd118;
  assign multm_reduce_mulb1_cq118 = xn2 & multm_reduce_sd119;
  assign multm_reduce_mulb1_cq119 = xn2 & multm_reduce_sd120;
  assign multm_reduce_mulb1_cq120 = xn2 & multm_reduce_sd121;
  assign multm_reduce_mulb1_cq121 = xn2 & multm_reduce_sd122;
  assign multm_reduce_mulb1_cq122 = xn2 & multm_reduce_sd123;
  assign multm_reduce_mulb1_cq123 = xn2 & multm_reduce_sd124;
  assign multm_reduce_mulb1_cq124 = xn2 & multm_reduce_sd125;
  assign multm_reduce_mulb1_cq125 = xn2 & multm_reduce_sd126;
  assign multm_reduce_mulb1_cq126 = xn2 & multm_reduce_sd127;
  assign multm_reduce_mulb1_cq127 = xn2 & multm_reduce_sd128;
  assign multm_reduce_mulb1_cq128 = xn2 & multm_reduce_sd129;
  assign multm_reduce_mulb1_cq129 = xn2 & multm_reduce_sd130;
  assign multm_reduce_mulb1_cq130 = xn2 & multm_reduce_sd131;
  assign multm_reduce_mulb1_cq131 = xn2 & multm_reduce_sd132;
  assign multm_reduce_mulb1_cq132 = xn2 & multm_reduce_sd133;
  assign multm_reduce_mulb1_cq133 = xn2 & multm_reduce_sd134;
  assign multm_reduce_mulb1_cq134 = xn2 & multm_reduce_sd135;
  assign multm_reduce_mulb1_cq135 = xn2 & multm_reduce_sd136;
  assign multm_reduce_mulb1_cq136 = xn2 & multm_reduce_sd137;
  assign multm_reduce_mulb1_cq137 = xn2 & multm_reduce_sd138;
  assign multm_reduce_mulb1_cq138 = xn2 & multm_reduce_sd139;
  assign multm_reduce_mulb1_cq139 = xn2 & multm_reduce_sd140;
  assign multm_reduce_mulb1_cq140 = xn2 & multm_reduce_sd141;
  assign multm_reduce_mulb1_cq141 = xn2 & multm_reduce_sd142;
  assign multm_reduce_mulb1_cq142 = xn2 & multm_reduce_sd143;
  assign multm_reduce_mulb1_cq143 = xn2 & multm_reduce_sd144;
  assign multm_reduce_mulb1_cq144 = xn2 & multm_reduce_sd145;
  assign multm_reduce_mulb1_cq145 = xn2 & multm_reduce_sd146;
  assign multm_reduce_mulb1_cq146 = xn2 & multm_reduce_sd147;
  assign multm_reduce_mulb1_cq147 = xn2 & multm_reduce_sd148;
  assign multm_reduce_mulb1_cq148 = xn2 & multm_reduce_sd149;
  assign multm_reduce_mulb1_cq149 = xn2 & multm_reduce_sd150;
  assign multm_reduce_mulb1_cq150 = xn2 & multm_reduce_sd151;
  assign multm_reduce_mulb1_cq151 = xn2 & multm_reduce_sd152;
  assign multm_reduce_mulb1_cq152 = xn2 & multm_reduce_sd153;
  assign multm_reduce_mulb1_cq153 = xn2 & multm_reduce_sd154;
  assign multm_reduce_mulb1_cq154 = xn2 & multm_reduce_sd155;
  assign multm_reduce_mulb1_cq155 = xn2 & multm_reduce_sd156;
  assign multm_reduce_mulb1_cq156 = xn2 & multm_reduce_sd157;
  assign multm_reduce_mulb1_cq157 = xn2 & multm_reduce_sd158;
  assign multm_reduce_mulb1_cq158 = xn2 & multm_reduce_sd159;
  assign multm_reduce_mulb1_cq159 = xn2 & multm_reduce_sd160;
  assign multm_reduce_mulb1_cq160 = xn2 & multm_reduce_sd161;
  assign multm_reduce_mulb1_cq161 = xn2 & multm_reduce_sd162;
  assign multm_reduce_mulb1_cq162 = xn2 & multm_reduce_sd163;
  assign multm_reduce_mulb1_cq163 = xn2 & multm_reduce_sd164;
  assign multm_reduce_mulb1_cq164 = xn2 & multm_reduce_sd165;
  assign multm_reduce_mulb1_cq165 = xn2 & multm_reduce_sd166;
  assign multm_reduce_mulb1_cq166 = xn2 & multm_reduce_sd167;
  assign multm_reduce_mulb1_cq167 = xn2 & multm_reduce_sd168;
  assign multm_reduce_mulb1_cq168 = xn2 & multm_reduce_sd169;
  assign multm_reduce_mulb1_cq169 = xn2 & multm_reduce_sd170;
  assign multm_reduce_mulb1_cq170 = xn2 & multm_reduce_sd171;
  assign multm_reduce_mulb1_cq171 = xn2 & multm_reduce_sd172;
  assign multm_reduce_mulb1_cq172 = xn2 & multm_reduce_sd173;
  assign multm_reduce_mulb1_cq173 = xn2 & multm_reduce_sd174;
  assign multm_reduce_mulb1_cq174 = xn2 & multm_reduce_sd175;
  assign multm_reduce_mulb1_cq175 = xn2 & multm_reduce_sd176;
  assign multm_reduce_mulb1_cq176 = xn2 & multm_reduce_sd177;
  assign multm_reduce_mulb1_cq177 = xn2 & multm_reduce_sd178;
  assign multm_reduce_mulb1_cq178 = xn2 & multm_reduce_sd179;
  assign multm_reduce_mulb1_cq179 = xn2 & multm_reduce_sd180;
  assign multm_reduce_mulb1_cq180 = xn2 & multm_reduce_sd181;
  assign multm_reduce_mulb1_cq181 = xn2 & multm_reduce_sd182;
  assign multm_reduce_mulb1_cq182 = xn2 & multm_reduce_sd183;
  assign multm_reduce_mulb1_pc0 = multm_reduce_mulb1_sq0 & multm_reduce_qb2;
  assign multm_reduce_mulb1_pc1 = multm_reduce_mulb1_add3b_maj3b_or3b_wx0 | multm_reduce_mulb1_add3b_maj3b_xy0;
  assign multm_reduce_mulb1_pc2 = multm_reduce_mulb1_add3b_maj3b_or3b_wx1 | multm_reduce_mulb1_add3b_maj3b_xy1;
  assign multm_reduce_mulb1_pc3 = multm_reduce_mulb1_sq3 & multm_reduce_mulb1_cq2;
  assign multm_reduce_mulb1_pc4 = multm_reduce_mulb1_sq4 & multm_reduce_mulb1_cq3;
  assign multm_reduce_mulb1_pc5 = multm_reduce_mulb1_add3b_maj3b_or3b_wx4 | multm_reduce_mulb1_add3b_maj3b_xy4;
  assign multm_reduce_mulb1_pc6 = multm_reduce_mulb1_add3b_maj3b_or3b_wx5 | multm_reduce_mulb1_add3b_maj3b_xy5;
  assign multm_reduce_mulb1_pc7 = multm_reduce_mulb1_add3b_maj3b_or3b_wx6 | multm_reduce_mulb1_add3b_maj3b_xy6;
  assign multm_reduce_mulb1_pc8 = multm_reduce_mulb1_add3b_maj3b_or3b_wx7 | multm_reduce_mulb1_add3b_maj3b_xy7;
  assign multm_reduce_mulb1_pc9 = multm_reduce_mulb1_sq9 & multm_reduce_mulb1_cq8;
  assign multm_reduce_mulb1_pc10 = multm_reduce_mulb1_sq10 & multm_reduce_mulb1_cq9;
  assign multm_reduce_mulb1_pc11 = multm_reduce_mulb1_add3b_maj3b_or3b_wx10 | multm_reduce_mulb1_add3b_maj3b_xy10;
  assign multm_reduce_mulb1_pc12 = multm_reduce_mulb1_sq12 & multm_reduce_mulb1_cq11;
  assign multm_reduce_mulb1_pc13 = multm_reduce_mulb1_add3b_maj3b_or3b_wx12 | multm_reduce_mulb1_add3b_maj3b_xy12;
  assign multm_reduce_mulb1_pc14 = multm_reduce_mulb1_sq14 & multm_reduce_mulb1_cq13;
  assign multm_reduce_mulb1_pc15 = multm_reduce_mulb1_sq15 & multm_reduce_mulb1_cq14;
  assign multm_reduce_mulb1_pc16 = multm_reduce_mulb1_sq16 & multm_reduce_mulb1_cq15;
  assign multm_reduce_mulb1_pc17 = multm_reduce_mulb1_sq17 & multm_reduce_mulb1_cq16;
  assign multm_reduce_mulb1_pc18 = multm_reduce_mulb1_sq18 & multm_reduce_mulb1_cq17;
  assign multm_reduce_mulb1_pc19 = multm_reduce_mulb1_add3b_maj3b_or3b_wx18 | multm_reduce_mulb1_add3b_maj3b_xy18;
  assign multm_reduce_mulb1_pc20 = multm_reduce_mulb1_sq20 & multm_reduce_mulb1_cq19;
  assign multm_reduce_mulb1_pc21 = multm_reduce_mulb1_add3b_maj3b_or3b_wx20 | multm_reduce_mulb1_add3b_maj3b_xy20;
  assign multm_reduce_mulb1_pc22 = multm_reduce_mulb1_sq22 & multm_reduce_mulb1_cq21;
  assign multm_reduce_mulb1_pc23 = multm_reduce_mulb1_add3b_maj3b_or3b_wx22 | multm_reduce_mulb1_add3b_maj3b_xy22;
  assign multm_reduce_mulb1_pc24 = multm_reduce_mulb1_add3b_maj3b_or3b_wx23 | multm_reduce_mulb1_add3b_maj3b_xy23;
  assign multm_reduce_mulb1_pc25 = multm_reduce_mulb1_add3b_maj3b_or3b_wx24 | multm_reduce_mulb1_add3b_maj3b_xy24;
  assign multm_reduce_mulb1_pc26 = multm_reduce_mulb1_sq26 & multm_reduce_mulb1_cq25;
  assign multm_reduce_mulb1_pc27 = multm_reduce_mulb1_sq27 & multm_reduce_mulb1_cq26;
  assign multm_reduce_mulb1_pc28 = multm_reduce_mulb1_sq28 & multm_reduce_mulb1_cq27;
  assign multm_reduce_mulb1_pc29 = multm_reduce_mulb1_add3b_maj3b_or3b_wx28 | multm_reduce_mulb1_add3b_maj3b_xy28;
  assign multm_reduce_mulb1_pc30 = multm_reduce_mulb1_sq30 & multm_reduce_mulb1_cq29;
  assign multm_reduce_mulb1_pc31 = multm_reduce_mulb1_add3b_maj3b_or3b_wx30 | multm_reduce_mulb1_add3b_maj3b_xy30;
  assign multm_reduce_mulb1_pc32 = multm_reduce_mulb1_sq32 & multm_reduce_mulb1_cq31;
  assign multm_reduce_mulb1_pc33 = multm_reduce_mulb1_add3b_maj3b_or3b_wx32 | multm_reduce_mulb1_add3b_maj3b_xy32;
  assign multm_reduce_mulb1_pc34 = multm_reduce_mulb1_sq34 & multm_reduce_mulb1_cq33;
  assign multm_reduce_mulb1_pc35 = multm_reduce_mulb1_add3b_maj3b_or3b_wx34 | multm_reduce_mulb1_add3b_maj3b_xy34;
  assign multm_reduce_mulb1_pc36 = multm_reduce_mulb1_sq36 & multm_reduce_mulb1_cq35;
  assign multm_reduce_mulb1_pc37 = multm_reduce_mulb1_sq37 & multm_reduce_mulb1_cq36;
  assign multm_reduce_mulb1_pc38 = multm_reduce_mulb1_add3b_maj3b_or3b_wx37 | multm_reduce_mulb1_add3b_maj3b_xy37;
  assign multm_reduce_mulb1_pc39 = multm_reduce_mulb1_sq39 & multm_reduce_mulb1_cq38;
  assign multm_reduce_mulb1_pc40 = multm_reduce_mulb1_sq40 & multm_reduce_mulb1_cq39;
  assign multm_reduce_mulb1_pc41 = multm_reduce_mulb1_add3b_maj3b_or3b_wx40 | multm_reduce_mulb1_add3b_maj3b_xy40;
  assign multm_reduce_mulb1_pc42 = multm_reduce_mulb1_add3b_maj3b_or3b_wx41 | multm_reduce_mulb1_add3b_maj3b_xy41;
  assign multm_reduce_mulb1_pc43 = multm_reduce_mulb1_add3b_maj3b_or3b_wx42 | multm_reduce_mulb1_add3b_maj3b_xy42;
  assign multm_reduce_mulb1_pc44 = multm_reduce_mulb1_add3b_maj3b_or3b_wx43 | multm_reduce_mulb1_add3b_maj3b_xy43;
  assign multm_reduce_mulb1_pc45 = multm_reduce_mulb1_sq45 & multm_reduce_mulb1_cq44;
  assign multm_reduce_mulb1_pc46 = multm_reduce_mulb1_sq46 & multm_reduce_mulb1_cq45;
  assign multm_reduce_mulb1_pc47 = multm_reduce_mulb1_sq47 & multm_reduce_mulb1_cq46;
  assign multm_reduce_mulb1_pc48 = multm_reduce_mulb1_add3b_maj3b_or3b_wx47 | multm_reduce_mulb1_add3b_maj3b_xy47;
  assign multm_reduce_mulb1_pc49 = multm_reduce_mulb1_add3b_maj3b_or3b_wx48 | multm_reduce_mulb1_add3b_maj3b_xy48;
  assign multm_reduce_mulb1_pc50 = multm_reduce_mulb1_sq50 & multm_reduce_mulb1_cq49;
  assign multm_reduce_mulb1_pc51 = multm_reduce_mulb1_sq51 & multm_reduce_mulb1_cq50;
  assign multm_reduce_mulb1_pc52 = multm_reduce_mulb1_add3b_maj3b_or3b_wx51 | multm_reduce_mulb1_add3b_maj3b_xy51;
  assign multm_reduce_mulb1_pc53 = multm_reduce_mulb1_add3b_maj3b_or3b_wx52 | multm_reduce_mulb1_add3b_maj3b_xy52;
  assign multm_reduce_mulb1_pc54 = multm_reduce_mulb1_add3b_maj3b_or3b_wx53 | multm_reduce_mulb1_add3b_maj3b_xy53;
  assign multm_reduce_mulb1_pc55 = multm_reduce_mulb1_add3b_maj3b_or3b_wx54 | multm_reduce_mulb1_add3b_maj3b_xy54;
  assign multm_reduce_mulb1_pc56 = multm_reduce_mulb1_add3b_maj3b_or3b_wx55 | multm_reduce_mulb1_add3b_maj3b_xy55;
  assign multm_reduce_mulb1_pc57 = multm_reduce_mulb1_sq57 & multm_reduce_mulb1_cq56;
  assign multm_reduce_mulb1_pc58 = multm_reduce_mulb1_add3b_maj3b_or3b_wx57 | multm_reduce_mulb1_add3b_maj3b_xy57;
  assign multm_reduce_mulb1_pc59 = multm_reduce_mulb1_sq59 & multm_reduce_mulb1_cq58;
  assign multm_reduce_mulb1_pc60 = multm_reduce_mulb1_sq60 & multm_reduce_mulb1_cq59;
  assign multm_reduce_mulb1_pc61 = multm_reduce_mulb1_sq61 & multm_reduce_mulb1_cq60;
  assign multm_reduce_mulb1_pc62 = multm_reduce_mulb1_sq62 & multm_reduce_mulb1_cq61;
  assign multm_reduce_mulb1_pc63 = multm_reduce_mulb1_add3b_maj3b_or3b_wx62 | multm_reduce_mulb1_add3b_maj3b_xy62;
  assign multm_reduce_mulb1_pc64 = multm_reduce_mulb1_sq64 & multm_reduce_mulb1_cq63;
  assign multm_reduce_mulb1_pc65 = multm_reduce_mulb1_sq65 & multm_reduce_mulb1_cq64;
  assign multm_reduce_mulb1_pc66 = multm_reduce_mulb1_sq66 & multm_reduce_mulb1_cq65;
  assign multm_reduce_mulb1_pc67 = multm_reduce_mulb1_add3b_maj3b_or3b_wx66 | multm_reduce_mulb1_add3b_maj3b_xy66;
  assign multm_reduce_mulb1_pc68 = multm_reduce_mulb1_sq68 & multm_reduce_mulb1_cq67;
  assign multm_reduce_mulb1_pc69 = multm_reduce_mulb1_add3b_maj3b_or3b_wx68 | multm_reduce_mulb1_add3b_maj3b_xy68;
  assign multm_reduce_mulb1_pc70 = multm_reduce_mulb1_add3b_maj3b_or3b_wx69 | multm_reduce_mulb1_add3b_maj3b_xy69;
  assign multm_reduce_mulb1_pc71 = multm_reduce_mulb1_sq71 & multm_reduce_mulb1_cq70;
  assign multm_reduce_mulb1_pc72 = multm_reduce_mulb1_add3b_maj3b_or3b_wx71 | multm_reduce_mulb1_add3b_maj3b_xy71;
  assign multm_reduce_mulb1_pc73 = multm_reduce_mulb1_sq73 & multm_reduce_mulb1_cq72;
  assign multm_reduce_mulb1_pc74 = multm_reduce_mulb1_add3b_maj3b_or3b_wx73 | multm_reduce_mulb1_add3b_maj3b_xy73;
  assign multm_reduce_mulb1_pc75 = multm_reduce_mulb1_add3b_maj3b_or3b_wx74 | multm_reduce_mulb1_add3b_maj3b_xy74;
  assign multm_reduce_mulb1_pc76 = multm_reduce_mulb1_sq76 & multm_reduce_mulb1_cq75;
  assign multm_reduce_mulb1_pc77 = multm_reduce_mulb1_sq77 & multm_reduce_mulb1_cq76;
  assign multm_reduce_mulb1_pc78 = multm_reduce_mulb1_sq78 & multm_reduce_mulb1_cq77;
  assign multm_reduce_mulb1_pc79 = multm_reduce_mulb1_sq79 & multm_reduce_mulb1_cq78;
  assign multm_reduce_mulb1_pc80 = multm_reduce_mulb1_add3b_maj3b_or3b_wx79 | multm_reduce_mulb1_add3b_maj3b_xy79;
  assign multm_reduce_mulb1_pc81 = multm_reduce_mulb1_add3b_maj3b_or3b_wx80 | multm_reduce_mulb1_add3b_maj3b_xy80;
  assign multm_reduce_mulb1_pc82 = multm_reduce_mulb1_sq82 & multm_reduce_mulb1_cq81;
  assign multm_reduce_mulb1_pc83 = multm_reduce_mulb1_add3b_maj3b_or3b_wx82 | multm_reduce_mulb1_add3b_maj3b_xy82;
  assign multm_reduce_mulb1_pc84 = multm_reduce_mulb1_sq84 & multm_reduce_mulb1_cq83;
  assign multm_reduce_mulb1_pc85 = multm_reduce_mulb1_sq85 & multm_reduce_mulb1_cq84;
  assign multm_reduce_mulb1_pc86 = multm_reduce_mulb1_sq86 & multm_reduce_mulb1_cq85;
  assign multm_reduce_mulb1_pc87 = multm_reduce_mulb1_add3b_maj3b_or3b_wx86 | multm_reduce_mulb1_add3b_maj3b_xy86;
  assign multm_reduce_mulb1_pc88 = multm_reduce_mulb1_sq88 & multm_reduce_mulb1_cq87;
  assign multm_reduce_mulb1_pc89 = multm_reduce_mulb1_add3b_maj3b_or3b_wx88 | multm_reduce_mulb1_add3b_maj3b_xy88;
  assign multm_reduce_mulb1_pc90 = multm_reduce_mulb1_sq90 & multm_reduce_mulb1_cq89;
  assign multm_reduce_mulb1_pc91 = multm_reduce_mulb1_add3b_maj3b_or3b_wx90 | multm_reduce_mulb1_add3b_maj3b_xy90;
  assign multm_reduce_mulb1_pc92 = multm_reduce_mulb1_add3b_maj3b_or3b_wx91 | multm_reduce_mulb1_add3b_maj3b_xy91;
  assign multm_reduce_mulb1_pc93 = multm_reduce_mulb1_sq93 & multm_reduce_mulb1_cq92;
  assign multm_reduce_mulb1_pc94 = multm_reduce_mulb1_sq94 & multm_reduce_mulb1_cq93;
  assign multm_reduce_mulb1_pc95 = multm_reduce_mulb1_sq95 & multm_reduce_mulb1_cq94;
  assign multm_reduce_mulb1_pc96 = multm_reduce_mulb1_sq96 & multm_reduce_mulb1_cq95;
  assign multm_reduce_mulb1_pc97 = multm_reduce_mulb1_add3b_maj3b_or3b_wx96 | multm_reduce_mulb1_add3b_maj3b_xy96;
  assign multm_reduce_mulb1_pc98 = multm_reduce_mulb1_sq98 & multm_reduce_mulb1_cq97;
  assign multm_reduce_mulb1_pc99 = multm_reduce_mulb1_sq99 & multm_reduce_mulb1_cq98;
  assign multm_reduce_mulb1_pc100 = multm_reduce_mulb1_add3b_maj3b_or3b_wx99 | multm_reduce_mulb1_add3b_maj3b_xy99;
  assign multm_reduce_mulb1_pc101 = multm_reduce_mulb1_add3b_maj3b_or3b_wx100 | multm_reduce_mulb1_add3b_maj3b_xy100;
  assign multm_reduce_mulb1_pc102 = multm_reduce_mulb1_add3b_maj3b_or3b_wx101 | multm_reduce_mulb1_add3b_maj3b_xy101;
  assign multm_reduce_mulb1_pc103 = multm_reduce_mulb1_add3b_maj3b_or3b_wx102 | multm_reduce_mulb1_add3b_maj3b_xy102;
  assign multm_reduce_mulb1_pc104 = multm_reduce_mulb1_sq104 & multm_reduce_mulb1_cq103;
  assign multm_reduce_mulb1_pc105 = multm_reduce_mulb1_add3b_maj3b_or3b_wx104 | multm_reduce_mulb1_add3b_maj3b_xy104;
  assign multm_reduce_mulb1_pc106 = multm_reduce_mulb1_add3b_maj3b_or3b_wx105 | multm_reduce_mulb1_add3b_maj3b_xy105;
  assign multm_reduce_mulb1_pc107 = multm_reduce_mulb1_sq107 & multm_reduce_mulb1_cq106;
  assign multm_reduce_mulb1_pc108 = multm_reduce_mulb1_add3b_maj3b_or3b_wx107 | multm_reduce_mulb1_add3b_maj3b_xy107;
  assign multm_reduce_mulb1_pc109 = multm_reduce_mulb1_add3b_maj3b_or3b_wx108 | multm_reduce_mulb1_add3b_maj3b_xy108;
  assign multm_reduce_mulb1_pc110 = multm_reduce_mulb1_add3b_maj3b_or3b_wx109 | multm_reduce_mulb1_add3b_maj3b_xy109;
  assign multm_reduce_mulb1_pc111 = multm_reduce_mulb1_add3b_maj3b_or3b_wx110 | multm_reduce_mulb1_add3b_maj3b_xy110;
  assign multm_reduce_mulb1_pc112 = multm_reduce_mulb1_sq112 & multm_reduce_mulb1_cq111;
  assign multm_reduce_mulb1_pc113 = multm_reduce_mulb1_add3b_maj3b_or3b_wx112 | multm_reduce_mulb1_add3b_maj3b_xy112;
  assign multm_reduce_mulb1_pc114 = multm_reduce_mulb1_sq114 & multm_reduce_mulb1_cq113;
  assign multm_reduce_mulb1_pc115 = multm_reduce_mulb1_add3b_maj3b_or3b_wx114 | multm_reduce_mulb1_add3b_maj3b_xy114;
  assign multm_reduce_mulb1_pc116 = multm_reduce_mulb1_sq116 & multm_reduce_mulb1_cq115;
  assign multm_reduce_mulb1_pc117 = multm_reduce_mulb1_sq117 & multm_reduce_mulb1_cq116;
  assign multm_reduce_mulb1_pc118 = multm_reduce_mulb1_add3b_maj3b_or3b_wx117 | multm_reduce_mulb1_add3b_maj3b_xy117;
  assign multm_reduce_mulb1_pc119 = multm_reduce_mulb1_add3b_maj3b_or3b_wx118 | multm_reduce_mulb1_add3b_maj3b_xy118;
  assign multm_reduce_mulb1_pc120 = multm_reduce_mulb1_add3b_maj3b_or3b_wx119 | multm_reduce_mulb1_add3b_maj3b_xy119;
  assign multm_reduce_mulb1_pc121 = multm_reduce_mulb1_add3b_maj3b_or3b_wx120 | multm_reduce_mulb1_add3b_maj3b_xy120;
  assign multm_reduce_mulb1_pc122 = multm_reduce_mulb1_add3b_maj3b_or3b_wx121 | multm_reduce_mulb1_add3b_maj3b_xy121;
  assign multm_reduce_mulb1_pc123 = multm_reduce_mulb1_add3b_maj3b_or3b_wx122 | multm_reduce_mulb1_add3b_maj3b_xy122;
  assign multm_reduce_mulb1_pc124 = multm_reduce_mulb1_add3b_maj3b_or3b_wx123 | multm_reduce_mulb1_add3b_maj3b_xy123;
  assign multm_reduce_mulb1_pc125 = multm_reduce_mulb1_sq125 & multm_reduce_mulb1_cq124;
  assign multm_reduce_mulb1_pc126 = multm_reduce_mulb1_sq126 & multm_reduce_mulb1_cq125;
  assign multm_reduce_mulb1_pc127 = multm_reduce_mulb1_sq127 & multm_reduce_mulb1_cq126;
  assign multm_reduce_mulb1_pc128 = multm_reduce_mulb1_sq128 & multm_reduce_mulb1_cq127;
  assign multm_reduce_mulb1_pc129 = multm_reduce_mulb1_add3b_maj3b_or3b_wx128 | multm_reduce_mulb1_add3b_maj3b_xy128;
  assign multm_reduce_mulb1_pc130 = multm_reduce_mulb1_sq130 & multm_reduce_mulb1_cq129;
  assign multm_reduce_mulb1_pc131 = multm_reduce_mulb1_add3b_maj3b_or3b_wx130 | multm_reduce_mulb1_add3b_maj3b_xy130;
  assign multm_reduce_mulb1_pc132 = multm_reduce_mulb1_sq132 & multm_reduce_mulb1_cq131;
  assign multm_reduce_mulb1_pc133 = multm_reduce_mulb1_add3b_maj3b_or3b_wx132 | multm_reduce_mulb1_add3b_maj3b_xy132;
  assign multm_reduce_mulb1_pc134 = multm_reduce_mulb1_sq134 & multm_reduce_mulb1_cq133;
  assign multm_reduce_mulb1_pc135 = multm_reduce_mulb1_sq135 & multm_reduce_mulb1_cq134;
  assign multm_reduce_mulb1_pc136 = multm_reduce_mulb1_add3b_maj3b_or3b_wx135 | multm_reduce_mulb1_add3b_maj3b_xy135;
  assign multm_reduce_mulb1_pc137 = multm_reduce_mulb1_add3b_maj3b_or3b_wx136 | multm_reduce_mulb1_add3b_maj3b_xy136;
  assign multm_reduce_mulb1_pc138 = multm_reduce_mulb1_sq138 & multm_reduce_mulb1_cq137;
  assign multm_reduce_mulb1_pc139 = multm_reduce_mulb1_sq139 & multm_reduce_mulb1_cq138;
  assign multm_reduce_mulb1_pc140 = multm_reduce_mulb1_sq140 & multm_reduce_mulb1_cq139;
  assign multm_reduce_mulb1_pc141 = multm_reduce_mulb1_add3b_maj3b_or3b_wx140 | multm_reduce_mulb1_add3b_maj3b_xy140;
  assign multm_reduce_mulb1_pc142 = multm_reduce_mulb1_add3b_maj3b_or3b_wx141 | multm_reduce_mulb1_add3b_maj3b_xy141;
  assign multm_reduce_mulb1_pc143 = multm_reduce_mulb1_add3b_maj3b_or3b_wx142 | multm_reduce_mulb1_add3b_maj3b_xy142;
  assign multm_reduce_mulb1_pc144 = multm_reduce_mulb1_add3b_maj3b_or3b_wx143 | multm_reduce_mulb1_add3b_maj3b_xy143;
  assign multm_reduce_mulb1_pc145 = multm_reduce_mulb1_add3b_maj3b_or3b_wx144 | multm_reduce_mulb1_add3b_maj3b_xy144;
  assign multm_reduce_mulb1_pc146 = multm_reduce_mulb1_sq146 & multm_reduce_mulb1_cq145;
  assign multm_reduce_mulb1_pc147 = multm_reduce_mulb1_sq147 & multm_reduce_mulb1_cq146;
  assign multm_reduce_mulb1_pc148 = multm_reduce_mulb1_add3b_maj3b_or3b_wx147 | multm_reduce_mulb1_add3b_maj3b_xy147;
  assign multm_reduce_mulb1_pc149 = multm_reduce_mulb1_sq149 & multm_reduce_mulb1_cq148;
  assign multm_reduce_mulb1_pc150 = multm_reduce_mulb1_sq150 & multm_reduce_mulb1_cq149;
  assign multm_reduce_mulb1_pc151 = multm_reduce_mulb1_add3b_maj3b_or3b_wx150 | multm_reduce_mulb1_add3b_maj3b_xy150;
  assign multm_reduce_mulb1_pc152 = multm_reduce_mulb1_add3b_maj3b_or3b_wx151 | multm_reduce_mulb1_add3b_maj3b_xy151;
  assign multm_reduce_mulb1_pc153 = multm_reduce_mulb1_add3b_maj3b_or3b_wx152 | multm_reduce_mulb1_add3b_maj3b_xy152;
  assign multm_reduce_mulb1_pc154 = multm_reduce_mulb1_add3b_maj3b_or3b_wx153 | multm_reduce_mulb1_add3b_maj3b_xy153;
  assign multm_reduce_mulb1_pc155 = multm_reduce_mulb1_sq155 & multm_reduce_mulb1_cq154;
  assign multm_reduce_mulb1_pc156 = multm_reduce_mulb1_add3b_maj3b_or3b_wx155 | multm_reduce_mulb1_add3b_maj3b_xy155;
  assign multm_reduce_mulb1_pc157 = multm_reduce_mulb1_add3b_maj3b_or3b_wx156 | multm_reduce_mulb1_add3b_maj3b_xy156;
  assign multm_reduce_mulb1_pc158 = multm_reduce_mulb1_add3b_maj3b_or3b_wx157 | multm_reduce_mulb1_add3b_maj3b_xy157;
  assign multm_reduce_mulb1_pc159 = multm_reduce_mulb1_add3b_maj3b_or3b_wx158 | multm_reduce_mulb1_add3b_maj3b_xy158;
  assign multm_reduce_mulb1_pc160 = multm_reduce_mulb1_add3b_maj3b_or3b_wx159 | multm_reduce_mulb1_add3b_maj3b_xy159;
  assign multm_reduce_mulb1_pc161 = multm_reduce_mulb1_add3b_maj3b_or3b_wx160 | multm_reduce_mulb1_add3b_maj3b_xy160;
  assign multm_reduce_mulb1_pc162 = multm_reduce_mulb1_sq162 & multm_reduce_mulb1_cq161;
  assign multm_reduce_mulb1_pc163 = multm_reduce_mulb1_add3b_maj3b_or3b_wx162 | multm_reduce_mulb1_add3b_maj3b_xy162;
  assign multm_reduce_mulb1_pc164 = multm_reduce_mulb1_sq164 & multm_reduce_mulb1_cq163;
  assign multm_reduce_mulb1_pc165 = multm_reduce_mulb1_sq165 & multm_reduce_mulb1_cq164;
  assign multm_reduce_mulb1_pc166 = multm_reduce_mulb1_sq166 & multm_reduce_mulb1_cq165;
  assign multm_reduce_mulb1_pc167 = multm_reduce_mulb1_add3b_maj3b_or3b_wx166 | multm_reduce_mulb1_add3b_maj3b_xy166;
  assign multm_reduce_mulb1_pc168 = multm_reduce_mulb1_sq168 & multm_reduce_mulb1_cq167;
  assign multm_reduce_mulb1_pc169 = multm_reduce_mulb1_sq169 & multm_reduce_mulb1_cq168;
  assign multm_reduce_mulb1_pc170 = multm_reduce_mulb1_sq170 & multm_reduce_mulb1_cq169;
  assign multm_reduce_mulb1_pc171 = multm_reduce_mulb1_sq171 & multm_reduce_mulb1_cq170;
  assign multm_reduce_mulb1_pc172 = multm_reduce_mulb1_add3b_maj3b_or3b_wx171 | multm_reduce_mulb1_add3b_maj3b_xy171;
  assign multm_reduce_mulb1_pc173 = multm_reduce_mulb1_add3b_maj3b_or3b_wx172 | multm_reduce_mulb1_add3b_maj3b_xy172;
  assign multm_reduce_mulb1_pc174 = multm_reduce_mulb1_add3b_maj3b_or3b_wx173 | multm_reduce_mulb1_add3b_maj3b_xy173;
  assign multm_reduce_mulb1_pc175 = multm_reduce_mulb1_add3b_maj3b_or3b_wx174 | multm_reduce_mulb1_add3b_maj3b_xy174;
  assign multm_reduce_mulb1_pc176 = multm_reduce_mulb1_add3b_maj3b_or3b_wx175 | multm_reduce_mulb1_add3b_maj3b_xy175;
  assign multm_reduce_mulb1_pc177 = multm_reduce_mulb1_sq177 & multm_reduce_mulb1_cq176;
  assign multm_reduce_mulb1_pc178 = multm_reduce_mulb1_sq178 & multm_reduce_mulb1_cq177;
  assign multm_reduce_mulb1_pc179 = multm_reduce_mulb1_sq179 & multm_reduce_mulb1_cq178;
  assign multm_reduce_mulb1_pc180 = multm_reduce_mulb1_add3b_maj3b_or3b_wx179 | multm_reduce_mulb1_add3b_maj3b_xy179;
  assign multm_reduce_mulb1_pc181 = multm_reduce_mulb1_sq181 & multm_reduce_mulb1_cq180;
  assign multm_reduce_mulb1_pc182 = multm_reduce_mulb1_add3b_maj3b_or3b_wx181 | multm_reduce_mulb1_add3b_maj3b_xy181;
  assign multm_reduce_mulb1_ps0 = multm_reduce_mulb1_add3b_xor3b_wx0 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps1 = multm_reduce_mulb1_add3b_xor3b_wx1 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps2 = multm_reduce_mulb1_sq3 ^ multm_reduce_mulb1_cq2;
  assign multm_reduce_mulb1_ps3 = multm_reduce_mulb1_sq4 ^ multm_reduce_mulb1_cq3;
  assign multm_reduce_mulb1_ps4 = multm_reduce_mulb1_add3b_xor3b_wx4 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps5 = multm_reduce_mulb1_add3b_xor3b_wx5 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps6 = multm_reduce_mulb1_add3b_xor3b_wx6 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps7 = multm_reduce_mulb1_add3b_xor3b_wx7 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps8 = multm_reduce_mulb1_sq9 ^ multm_reduce_mulb1_cq8;
  assign multm_reduce_mulb1_ps9 = multm_reduce_mulb1_sq10 ^ multm_reduce_mulb1_cq9;
  assign multm_reduce_mulb1_ps10 = multm_reduce_mulb1_add3b_xor3b_wx10 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps11 = multm_reduce_mulb1_sq12 ^ multm_reduce_mulb1_cq11;
  assign multm_reduce_mulb1_ps12 = multm_reduce_mulb1_add3b_xor3b_wx12 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps13 = multm_reduce_mulb1_sq14 ^ multm_reduce_mulb1_cq13;
  assign multm_reduce_mulb1_ps14 = multm_reduce_mulb1_sq15 ^ multm_reduce_mulb1_cq14;
  assign multm_reduce_mulb1_ps15 = multm_reduce_mulb1_sq16 ^ multm_reduce_mulb1_cq15;
  assign multm_reduce_mulb1_ps16 = multm_reduce_mulb1_sq17 ^ multm_reduce_mulb1_cq16;
  assign multm_reduce_mulb1_ps17 = multm_reduce_mulb1_sq18 ^ multm_reduce_mulb1_cq17;
  assign multm_reduce_mulb1_ps18 = multm_reduce_mulb1_add3b_xor3b_wx18 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps19 = multm_reduce_mulb1_sq20 ^ multm_reduce_mulb1_cq19;
  assign multm_reduce_mulb1_ps20 = multm_reduce_mulb1_add3b_xor3b_wx20 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps21 = multm_reduce_mulb1_sq22 ^ multm_reduce_mulb1_cq21;
  assign multm_reduce_mulb1_ps22 = multm_reduce_mulb1_add3b_xor3b_wx22 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps23 = multm_reduce_mulb1_add3b_xor3b_wx23 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps24 = multm_reduce_mulb1_add3b_xor3b_wx24 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps25 = multm_reduce_mulb1_sq26 ^ multm_reduce_mulb1_cq25;
  assign multm_reduce_mulb1_ps26 = multm_reduce_mulb1_sq27 ^ multm_reduce_mulb1_cq26;
  assign multm_reduce_mulb1_ps27 = multm_reduce_mulb1_sq28 ^ multm_reduce_mulb1_cq27;
  assign multm_reduce_mulb1_ps28 = multm_reduce_mulb1_add3b_xor3b_wx28 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps29 = multm_reduce_mulb1_sq30 ^ multm_reduce_mulb1_cq29;
  assign multm_reduce_mulb1_ps30 = multm_reduce_mulb1_add3b_xor3b_wx30 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps31 = multm_reduce_mulb1_sq32 ^ multm_reduce_mulb1_cq31;
  assign multm_reduce_mulb1_ps32 = multm_reduce_mulb1_add3b_xor3b_wx32 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps33 = multm_reduce_mulb1_sq34 ^ multm_reduce_mulb1_cq33;
  assign multm_reduce_mulb1_ps34 = multm_reduce_mulb1_add3b_xor3b_wx34 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps35 = multm_reduce_mulb1_sq36 ^ multm_reduce_mulb1_cq35;
  assign multm_reduce_mulb1_ps36 = multm_reduce_mulb1_sq37 ^ multm_reduce_mulb1_cq36;
  assign multm_reduce_mulb1_ps37 = multm_reduce_mulb1_add3b_xor3b_wx37 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps38 = multm_reduce_mulb1_sq39 ^ multm_reduce_mulb1_cq38;
  assign multm_reduce_mulb1_ps39 = multm_reduce_mulb1_sq40 ^ multm_reduce_mulb1_cq39;
  assign multm_reduce_mulb1_ps40 = multm_reduce_mulb1_add3b_xor3b_wx40 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps41 = multm_reduce_mulb1_add3b_xor3b_wx41 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps42 = multm_reduce_mulb1_add3b_xor3b_wx42 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps43 = multm_reduce_mulb1_add3b_xor3b_wx43 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps44 = multm_reduce_mulb1_sq45 ^ multm_reduce_mulb1_cq44;
  assign multm_reduce_mulb1_ps45 = multm_reduce_mulb1_sq46 ^ multm_reduce_mulb1_cq45;
  assign multm_reduce_mulb1_ps46 = multm_reduce_mulb1_sq47 ^ multm_reduce_mulb1_cq46;
  assign multm_reduce_mulb1_ps47 = multm_reduce_mulb1_add3b_xor3b_wx47 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps48 = multm_reduce_mulb1_add3b_xor3b_wx48 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps49 = multm_reduce_mulb1_sq50 ^ multm_reduce_mulb1_cq49;
  assign multm_reduce_mulb1_ps50 = multm_reduce_mulb1_sq51 ^ multm_reduce_mulb1_cq50;
  assign multm_reduce_mulb1_ps51 = multm_reduce_mulb1_add3b_xor3b_wx51 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps52 = multm_reduce_mulb1_add3b_xor3b_wx52 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps53 = multm_reduce_mulb1_add3b_xor3b_wx53 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps54 = multm_reduce_mulb1_add3b_xor3b_wx54 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps55 = multm_reduce_mulb1_add3b_xor3b_wx55 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps56 = multm_reduce_mulb1_sq57 ^ multm_reduce_mulb1_cq56;
  assign multm_reduce_mulb1_ps57 = multm_reduce_mulb1_add3b_xor3b_wx57 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps58 = multm_reduce_mulb1_sq59 ^ multm_reduce_mulb1_cq58;
  assign multm_reduce_mulb1_ps59 = multm_reduce_mulb1_sq60 ^ multm_reduce_mulb1_cq59;
  assign multm_reduce_mulb1_ps60 = multm_reduce_mulb1_sq61 ^ multm_reduce_mulb1_cq60;
  assign multm_reduce_mulb1_ps61 = multm_reduce_mulb1_sq62 ^ multm_reduce_mulb1_cq61;
  assign multm_reduce_mulb1_ps62 = multm_reduce_mulb1_add3b_xor3b_wx62 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps63 = multm_reduce_mulb1_sq64 ^ multm_reduce_mulb1_cq63;
  assign multm_reduce_mulb1_ps64 = multm_reduce_mulb1_sq65 ^ multm_reduce_mulb1_cq64;
  assign multm_reduce_mulb1_ps65 = multm_reduce_mulb1_sq66 ^ multm_reduce_mulb1_cq65;
  assign multm_reduce_mulb1_ps66 = multm_reduce_mulb1_add3b_xor3b_wx66 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps67 = multm_reduce_mulb1_sq68 ^ multm_reduce_mulb1_cq67;
  assign multm_reduce_mulb1_ps68 = multm_reduce_mulb1_add3b_xor3b_wx68 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps69 = multm_reduce_mulb1_add3b_xor3b_wx69 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps70 = multm_reduce_mulb1_sq71 ^ multm_reduce_mulb1_cq70;
  assign multm_reduce_mulb1_ps71 = multm_reduce_mulb1_add3b_xor3b_wx71 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps72 = multm_reduce_mulb1_sq73 ^ multm_reduce_mulb1_cq72;
  assign multm_reduce_mulb1_ps73 = multm_reduce_mulb1_add3b_xor3b_wx73 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps74 = multm_reduce_mulb1_add3b_xor3b_wx74 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps75 = multm_reduce_mulb1_sq76 ^ multm_reduce_mulb1_cq75;
  assign multm_reduce_mulb1_ps76 = multm_reduce_mulb1_sq77 ^ multm_reduce_mulb1_cq76;
  assign multm_reduce_mulb1_ps77 = multm_reduce_mulb1_sq78 ^ multm_reduce_mulb1_cq77;
  assign multm_reduce_mulb1_ps78 = multm_reduce_mulb1_sq79 ^ multm_reduce_mulb1_cq78;
  assign multm_reduce_mulb1_ps79 = multm_reduce_mulb1_add3b_xor3b_wx79 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps80 = multm_reduce_mulb1_add3b_xor3b_wx80 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps81 = multm_reduce_mulb1_sq82 ^ multm_reduce_mulb1_cq81;
  assign multm_reduce_mulb1_ps82 = multm_reduce_mulb1_add3b_xor3b_wx82 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps83 = multm_reduce_mulb1_sq84 ^ multm_reduce_mulb1_cq83;
  assign multm_reduce_mulb1_ps84 = multm_reduce_mulb1_sq85 ^ multm_reduce_mulb1_cq84;
  assign multm_reduce_mulb1_ps85 = multm_reduce_mulb1_sq86 ^ multm_reduce_mulb1_cq85;
  assign multm_reduce_mulb1_ps86 = multm_reduce_mulb1_add3b_xor3b_wx86 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps87 = multm_reduce_mulb1_sq88 ^ multm_reduce_mulb1_cq87;
  assign multm_reduce_mulb1_ps88 = multm_reduce_mulb1_add3b_xor3b_wx88 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps89 = multm_reduce_mulb1_sq90 ^ multm_reduce_mulb1_cq89;
  assign multm_reduce_mulb1_ps90 = multm_reduce_mulb1_add3b_xor3b_wx90 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps91 = multm_reduce_mulb1_add3b_xor3b_wx91 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps92 = multm_reduce_mulb1_sq93 ^ multm_reduce_mulb1_cq92;
  assign multm_reduce_mulb1_ps93 = multm_reduce_mulb1_sq94 ^ multm_reduce_mulb1_cq93;
  assign multm_reduce_mulb1_ps94 = multm_reduce_mulb1_sq95 ^ multm_reduce_mulb1_cq94;
  assign multm_reduce_mulb1_ps95 = multm_reduce_mulb1_sq96 ^ multm_reduce_mulb1_cq95;
  assign multm_reduce_mulb1_ps96 = multm_reduce_mulb1_add3b_xor3b_wx96 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps97 = multm_reduce_mulb1_sq98 ^ multm_reduce_mulb1_cq97;
  assign multm_reduce_mulb1_ps98 = multm_reduce_mulb1_sq99 ^ multm_reduce_mulb1_cq98;
  assign multm_reduce_mulb1_ps99 = multm_reduce_mulb1_add3b_xor3b_wx99 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps100 = multm_reduce_mulb1_add3b_xor3b_wx100 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps101 = multm_reduce_mulb1_add3b_xor3b_wx101 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps102 = multm_reduce_mulb1_add3b_xor3b_wx102 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps103 = multm_reduce_mulb1_sq104 ^ multm_reduce_mulb1_cq103;
  assign multm_reduce_mulb1_ps104 = multm_reduce_mulb1_add3b_xor3b_wx104 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps105 = multm_reduce_mulb1_add3b_xor3b_wx105 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps106 = multm_reduce_mulb1_sq107 ^ multm_reduce_mulb1_cq106;
  assign multm_reduce_mulb1_ps107 = multm_reduce_mulb1_add3b_xor3b_wx107 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps108 = multm_reduce_mulb1_add3b_xor3b_wx108 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps109 = multm_reduce_mulb1_add3b_xor3b_wx109 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps110 = multm_reduce_mulb1_add3b_xor3b_wx110 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps111 = multm_reduce_mulb1_sq112 ^ multm_reduce_mulb1_cq111;
  assign multm_reduce_mulb1_ps112 = multm_reduce_mulb1_add3b_xor3b_wx112 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps113 = multm_reduce_mulb1_sq114 ^ multm_reduce_mulb1_cq113;
  assign multm_reduce_mulb1_ps114 = multm_reduce_mulb1_add3b_xor3b_wx114 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps115 = multm_reduce_mulb1_sq116 ^ multm_reduce_mulb1_cq115;
  assign multm_reduce_mulb1_ps116 = multm_reduce_mulb1_sq117 ^ multm_reduce_mulb1_cq116;
  assign multm_reduce_mulb1_ps117 = multm_reduce_mulb1_add3b_xor3b_wx117 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps118 = multm_reduce_mulb1_add3b_xor3b_wx118 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps119 = multm_reduce_mulb1_add3b_xor3b_wx119 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps120 = multm_reduce_mulb1_add3b_xor3b_wx120 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps121 = multm_reduce_mulb1_add3b_xor3b_wx121 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps122 = multm_reduce_mulb1_add3b_xor3b_wx122 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps123 = multm_reduce_mulb1_add3b_xor3b_wx123 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps124 = multm_reduce_mulb1_sq125 ^ multm_reduce_mulb1_cq124;
  assign multm_reduce_mulb1_ps125 = multm_reduce_mulb1_sq126 ^ multm_reduce_mulb1_cq125;
  assign multm_reduce_mulb1_ps126 = multm_reduce_mulb1_sq127 ^ multm_reduce_mulb1_cq126;
  assign multm_reduce_mulb1_ps127 = multm_reduce_mulb1_sq128 ^ multm_reduce_mulb1_cq127;
  assign multm_reduce_mulb1_ps128 = multm_reduce_mulb1_add3b_xor3b_wx128 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps129 = multm_reduce_mulb1_sq130 ^ multm_reduce_mulb1_cq129;
  assign multm_reduce_mulb1_ps130 = multm_reduce_mulb1_add3b_xor3b_wx130 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps131 = multm_reduce_mulb1_sq132 ^ multm_reduce_mulb1_cq131;
  assign multm_reduce_mulb1_ps132 = multm_reduce_mulb1_add3b_xor3b_wx132 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps133 = multm_reduce_mulb1_sq134 ^ multm_reduce_mulb1_cq133;
  assign multm_reduce_mulb1_ps134 = multm_reduce_mulb1_sq135 ^ multm_reduce_mulb1_cq134;
  assign multm_reduce_mulb1_ps135 = multm_reduce_mulb1_add3b_xor3b_wx135 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps136 = multm_reduce_mulb1_add3b_xor3b_wx136 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps137 = multm_reduce_mulb1_sq138 ^ multm_reduce_mulb1_cq137;
  assign multm_reduce_mulb1_ps138 = multm_reduce_mulb1_sq139 ^ multm_reduce_mulb1_cq138;
  assign multm_reduce_mulb1_ps139 = multm_reduce_mulb1_sq140 ^ multm_reduce_mulb1_cq139;
  assign multm_reduce_mulb1_ps140 = multm_reduce_mulb1_add3b_xor3b_wx140 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps141 = multm_reduce_mulb1_add3b_xor3b_wx141 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps142 = multm_reduce_mulb1_add3b_xor3b_wx142 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps143 = multm_reduce_mulb1_add3b_xor3b_wx143 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps144 = multm_reduce_mulb1_add3b_xor3b_wx144 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps145 = multm_reduce_mulb1_sq146 ^ multm_reduce_mulb1_cq145;
  assign multm_reduce_mulb1_ps146 = multm_reduce_mulb1_sq147 ^ multm_reduce_mulb1_cq146;
  assign multm_reduce_mulb1_ps147 = multm_reduce_mulb1_add3b_xor3b_wx147 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps148 = multm_reduce_mulb1_sq149 ^ multm_reduce_mulb1_cq148;
  assign multm_reduce_mulb1_ps149 = multm_reduce_mulb1_sq150 ^ multm_reduce_mulb1_cq149;
  assign multm_reduce_mulb1_ps150 = multm_reduce_mulb1_add3b_xor3b_wx150 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps151 = multm_reduce_mulb1_add3b_xor3b_wx151 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps152 = multm_reduce_mulb1_add3b_xor3b_wx152 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps153 = multm_reduce_mulb1_add3b_xor3b_wx153 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps154 = multm_reduce_mulb1_sq155 ^ multm_reduce_mulb1_cq154;
  assign multm_reduce_mulb1_ps155 = multm_reduce_mulb1_add3b_xor3b_wx155 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps156 = multm_reduce_mulb1_add3b_xor3b_wx156 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps157 = multm_reduce_mulb1_add3b_xor3b_wx157 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps158 = multm_reduce_mulb1_add3b_xor3b_wx158 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps159 = multm_reduce_mulb1_add3b_xor3b_wx159 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps160 = multm_reduce_mulb1_add3b_xor3b_wx160 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps161 = multm_reduce_mulb1_sq162 ^ multm_reduce_mulb1_cq161;
  assign multm_reduce_mulb1_ps162 = multm_reduce_mulb1_add3b_xor3b_wx162 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps163 = multm_reduce_mulb1_sq164 ^ multm_reduce_mulb1_cq163;
  assign multm_reduce_mulb1_ps164 = multm_reduce_mulb1_sq165 ^ multm_reduce_mulb1_cq164;
  assign multm_reduce_mulb1_ps165 = multm_reduce_mulb1_sq166 ^ multm_reduce_mulb1_cq165;
  assign multm_reduce_mulb1_ps166 = multm_reduce_mulb1_add3b_xor3b_wx166 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps167 = multm_reduce_mulb1_sq168 ^ multm_reduce_mulb1_cq167;
  assign multm_reduce_mulb1_ps168 = multm_reduce_mulb1_sq169 ^ multm_reduce_mulb1_cq168;
  assign multm_reduce_mulb1_ps169 = multm_reduce_mulb1_sq170 ^ multm_reduce_mulb1_cq169;
  assign multm_reduce_mulb1_ps170 = multm_reduce_mulb1_sq171 ^ multm_reduce_mulb1_cq170;
  assign multm_reduce_mulb1_ps171 = multm_reduce_mulb1_add3b_xor3b_wx171 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps172 = multm_reduce_mulb1_add3b_xor3b_wx172 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps173 = multm_reduce_mulb1_add3b_xor3b_wx173 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps174 = multm_reduce_mulb1_add3b_xor3b_wx174 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps175 = multm_reduce_mulb1_add3b_xor3b_wx175 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps176 = multm_reduce_mulb1_sq177 ^ multm_reduce_mulb1_cq176;
  assign multm_reduce_mulb1_ps177 = multm_reduce_mulb1_sq178 ^ multm_reduce_mulb1_cq177;
  assign multm_reduce_mulb1_ps178 = multm_reduce_mulb1_sq179 ^ multm_reduce_mulb1_cq178;
  assign multm_reduce_mulb1_ps179 = multm_reduce_mulb1_add3b_xor3b_wx179 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_ps180 = multm_reduce_mulb1_sq181 ^ multm_reduce_mulb1_cq180;
  assign multm_reduce_mulb1_ps181 = multm_reduce_mulb1_add3b_xor3b_wx181 ^ multm_reduce_qb2;
  assign multm_reduce_mulb1_sq0 = xn2 & multm_reduce_sc0;
  assign multm_reduce_mulb1_sq1 = xn2 & multm_reduce_sc1;
  assign multm_reduce_mulb1_sq2 = xn2 & multm_reduce_sc2;
  assign multm_reduce_mulb1_sq3 = xn2 & multm_reduce_sc3;
  assign multm_reduce_mulb1_sq4 = xn2 & multm_reduce_sc4;
  assign multm_reduce_mulb1_sq5 = xn2 & multm_reduce_sc5;
  assign multm_reduce_mulb1_sq6 = xn2 & multm_reduce_sc6;
  assign multm_reduce_mulb1_sq7 = xn2 & multm_reduce_sc7;
  assign multm_reduce_mulb1_sq8 = xn2 & multm_reduce_sc8;
  assign multm_reduce_mulb1_sq9 = xn2 & multm_reduce_sc9;
  assign multm_reduce_mulb1_sq10 = xn2 & multm_reduce_sc10;
  assign multm_reduce_mulb1_sq11 = xn2 & multm_reduce_sc11;
  assign multm_reduce_mulb1_sq12 = xn2 & multm_reduce_sc12;
  assign multm_reduce_mulb1_sq13 = xn2 & multm_reduce_sc13;
  assign multm_reduce_mulb1_sq14 = xn2 & multm_reduce_sc14;
  assign multm_reduce_mulb1_sq15 = xn2 & multm_reduce_sc15;
  assign multm_reduce_mulb1_sq16 = xn2 & multm_reduce_sc16;
  assign multm_reduce_mulb1_sq17 = xn2 & multm_reduce_sc17;
  assign multm_reduce_mulb1_sq18 = xn2 & multm_reduce_sc18;
  assign multm_reduce_mulb1_sq19 = xn2 & multm_reduce_sc19;
  assign multm_reduce_mulb1_sq20 = xn2 & multm_reduce_sc20;
  assign multm_reduce_mulb1_sq21 = xn2 & multm_reduce_sc21;
  assign multm_reduce_mulb1_sq22 = xn2 & multm_reduce_sc22;
  assign multm_reduce_mulb1_sq23 = xn2 & multm_reduce_sc23;
  assign multm_reduce_mulb1_sq24 = xn2 & multm_reduce_sc24;
  assign multm_reduce_mulb1_sq25 = xn2 & multm_reduce_sc25;
  assign multm_reduce_mulb1_sq26 = xn2 & multm_reduce_sc26;
  assign multm_reduce_mulb1_sq27 = xn2 & multm_reduce_sc27;
  assign multm_reduce_mulb1_sq28 = xn2 & multm_reduce_sc28;
  assign multm_reduce_mulb1_sq29 = xn2 & multm_reduce_sc29;
  assign multm_reduce_mulb1_sq30 = xn2 & multm_reduce_sc30;
  assign multm_reduce_mulb1_sq31 = xn2 & multm_reduce_sc31;
  assign multm_reduce_mulb1_sq32 = xn2 & multm_reduce_sc32;
  assign multm_reduce_mulb1_sq33 = xn2 & multm_reduce_sc33;
  assign multm_reduce_mulb1_sq34 = xn2 & multm_reduce_sc34;
  assign multm_reduce_mulb1_sq35 = xn2 & multm_reduce_sc35;
  assign multm_reduce_mulb1_sq36 = xn2 & multm_reduce_sc36;
  assign multm_reduce_mulb1_sq37 = xn2 & multm_reduce_sc37;
  assign multm_reduce_mulb1_sq38 = xn2 & multm_reduce_sc38;
  assign multm_reduce_mulb1_sq39 = xn2 & multm_reduce_sc39;
  assign multm_reduce_mulb1_sq40 = xn2 & multm_reduce_sc40;
  assign multm_reduce_mulb1_sq41 = xn2 & multm_reduce_sc41;
  assign multm_reduce_mulb1_sq42 = xn2 & multm_reduce_sc42;
  assign multm_reduce_mulb1_sq43 = xn2 & multm_reduce_sc43;
  assign multm_reduce_mulb1_sq44 = xn2 & multm_reduce_sc44;
  assign multm_reduce_mulb1_sq45 = xn2 & multm_reduce_sc45;
  assign multm_reduce_mulb1_sq46 = xn2 & multm_reduce_sc46;
  assign multm_reduce_mulb1_sq47 = xn2 & multm_reduce_sc47;
  assign multm_reduce_mulb1_sq48 = xn2 & multm_reduce_sc48;
  assign multm_reduce_mulb1_sq49 = xn2 & multm_reduce_sc49;
  assign multm_reduce_mulb1_sq50 = xn2 & multm_reduce_sc50;
  assign multm_reduce_mulb1_sq51 = xn2 & multm_reduce_sc51;
  assign multm_reduce_mulb1_sq52 = xn2 & multm_reduce_sc52;
  assign multm_reduce_mulb1_sq53 = xn2 & multm_reduce_sc53;
  assign multm_reduce_mulb1_sq54 = xn2 & multm_reduce_sc54;
  assign multm_reduce_mulb1_sq55 = xn2 & multm_reduce_sc55;
  assign multm_reduce_mulb1_sq56 = xn2 & multm_reduce_sc56;
  assign multm_reduce_mulb1_sq57 = xn2 & multm_reduce_sc57;
  assign multm_reduce_mulb1_sq58 = xn2 & multm_reduce_sc58;
  assign multm_reduce_mulb1_sq59 = xn2 & multm_reduce_sc59;
  assign multm_reduce_mulb1_sq60 = xn2 & multm_reduce_sc60;
  assign multm_reduce_mulb1_sq61 = xn2 & multm_reduce_sc61;
  assign multm_reduce_mulb1_sq62 = xn2 & multm_reduce_sc62;
  assign multm_reduce_mulb1_sq63 = xn2 & multm_reduce_sc63;
  assign multm_reduce_mulb1_sq64 = xn2 & multm_reduce_sc64;
  assign multm_reduce_mulb1_sq65 = xn2 & multm_reduce_sc65;
  assign multm_reduce_mulb1_sq66 = xn2 & multm_reduce_sc66;
  assign multm_reduce_mulb1_sq67 = xn2 & multm_reduce_sc67;
  assign multm_reduce_mulb1_sq68 = xn2 & multm_reduce_sc68;
  assign multm_reduce_mulb1_sq69 = xn2 & multm_reduce_sc69;
  assign multm_reduce_mulb1_sq70 = xn2 & multm_reduce_sc70;
  assign multm_reduce_mulb1_sq71 = xn2 & multm_reduce_sc71;
  assign multm_reduce_mulb1_sq72 = xn2 & multm_reduce_sc72;
  assign multm_reduce_mulb1_sq73 = xn2 & multm_reduce_sc73;
  assign multm_reduce_mulb1_sq74 = xn2 & multm_reduce_sc74;
  assign multm_reduce_mulb1_sq75 = xn2 & multm_reduce_sc75;
  assign multm_reduce_mulb1_sq76 = xn2 & multm_reduce_sc76;
  assign multm_reduce_mulb1_sq77 = xn2 & multm_reduce_sc77;
  assign multm_reduce_mulb1_sq78 = xn2 & multm_reduce_sc78;
  assign multm_reduce_mulb1_sq79 = xn2 & multm_reduce_sc79;
  assign multm_reduce_mulb1_sq80 = xn2 & multm_reduce_sc80;
  assign multm_reduce_mulb1_sq81 = xn2 & multm_reduce_sc81;
  assign multm_reduce_mulb1_sq82 = xn2 & multm_reduce_sc82;
  assign multm_reduce_mulb1_sq83 = xn2 & multm_reduce_sc83;
  assign multm_reduce_mulb1_sq84 = xn2 & multm_reduce_sc84;
  assign multm_reduce_mulb1_sq85 = xn2 & multm_reduce_sc85;
  assign multm_reduce_mulb1_sq86 = xn2 & multm_reduce_sc86;
  assign multm_reduce_mulb1_sq87 = xn2 & multm_reduce_sc87;
  assign multm_reduce_mulb1_sq88 = xn2 & multm_reduce_sc88;
  assign multm_reduce_mulb1_sq89 = xn2 & multm_reduce_sc89;
  assign multm_reduce_mulb1_sq90 = xn2 & multm_reduce_sc90;
  assign multm_reduce_mulb1_sq91 = xn2 & multm_reduce_sc91;
  assign multm_reduce_mulb1_sq92 = xn2 & multm_reduce_sc92;
  assign multm_reduce_mulb1_sq93 = xn2 & multm_reduce_sc93;
  assign multm_reduce_mulb1_sq94 = xn2 & multm_reduce_sc94;
  assign multm_reduce_mulb1_sq95 = xn2 & multm_reduce_sc95;
  assign multm_reduce_mulb1_sq96 = xn2 & multm_reduce_sc96;
  assign multm_reduce_mulb1_sq97 = xn2 & multm_reduce_sc97;
  assign multm_reduce_mulb1_sq98 = xn2 & multm_reduce_sc98;
  assign multm_reduce_mulb1_sq99 = xn2 & multm_reduce_sc99;
  assign multm_reduce_mulb1_sq100 = xn2 & multm_reduce_sc100;
  assign multm_reduce_mulb1_sq101 = xn2 & multm_reduce_sc101;
  assign multm_reduce_mulb1_sq102 = xn2 & multm_reduce_sc102;
  assign multm_reduce_mulb1_sq103 = xn2 & multm_reduce_sc103;
  assign multm_reduce_mulb1_sq104 = xn2 & multm_reduce_sc104;
  assign multm_reduce_mulb1_sq105 = xn2 & multm_reduce_sc105;
  assign multm_reduce_mulb1_sq106 = xn2 & multm_reduce_sc106;
  assign multm_reduce_mulb1_sq107 = xn2 & multm_reduce_sc107;
  assign multm_reduce_mulb1_sq108 = xn2 & multm_reduce_sc108;
  assign multm_reduce_mulb1_sq109 = xn2 & multm_reduce_sc109;
  assign multm_reduce_mulb1_sq110 = xn2 & multm_reduce_sc110;
  assign multm_reduce_mulb1_sq111 = xn2 & multm_reduce_sc111;
  assign multm_reduce_mulb1_sq112 = xn2 & multm_reduce_sc112;
  assign multm_reduce_mulb1_sq113 = xn2 & multm_reduce_sc113;
  assign multm_reduce_mulb1_sq114 = xn2 & multm_reduce_sc114;
  assign multm_reduce_mulb1_sq115 = xn2 & multm_reduce_sc115;
  assign multm_reduce_mulb1_sq116 = xn2 & multm_reduce_sc116;
  assign multm_reduce_mulb1_sq117 = xn2 & multm_reduce_sc117;
  assign multm_reduce_mulb1_sq118 = xn2 & multm_reduce_sc118;
  assign multm_reduce_mulb1_sq119 = xn2 & multm_reduce_sc119;
  assign multm_reduce_mulb1_sq120 = xn2 & multm_reduce_sc120;
  assign multm_reduce_mulb1_sq121 = xn2 & multm_reduce_sc121;
  assign multm_reduce_mulb1_sq122 = xn2 & multm_reduce_sc122;
  assign multm_reduce_mulb1_sq123 = xn2 & multm_reduce_sc123;
  assign multm_reduce_mulb1_sq124 = xn2 & multm_reduce_sc124;
  assign multm_reduce_mulb1_sq125 = xn2 & multm_reduce_sc125;
  assign multm_reduce_mulb1_sq126 = xn2 & multm_reduce_sc126;
  assign multm_reduce_mulb1_sq127 = xn2 & multm_reduce_sc127;
  assign multm_reduce_mulb1_sq128 = xn2 & multm_reduce_sc128;
  assign multm_reduce_mulb1_sq129 = xn2 & multm_reduce_sc129;
  assign multm_reduce_mulb1_sq130 = xn2 & multm_reduce_sc130;
  assign multm_reduce_mulb1_sq131 = xn2 & multm_reduce_sc131;
  assign multm_reduce_mulb1_sq132 = xn2 & multm_reduce_sc132;
  assign multm_reduce_mulb1_sq133 = xn2 & multm_reduce_sc133;
  assign multm_reduce_mulb1_sq134 = xn2 & multm_reduce_sc134;
  assign multm_reduce_mulb1_sq135 = xn2 & multm_reduce_sc135;
  assign multm_reduce_mulb1_sq136 = xn2 & multm_reduce_sc136;
  assign multm_reduce_mulb1_sq137 = xn2 & multm_reduce_sc137;
  assign multm_reduce_mulb1_sq138 = xn2 & multm_reduce_sc138;
  assign multm_reduce_mulb1_sq139 = xn2 & multm_reduce_sc139;
  assign multm_reduce_mulb1_sq140 = xn2 & multm_reduce_sc140;
  assign multm_reduce_mulb1_sq141 = xn2 & multm_reduce_sc141;
  assign multm_reduce_mulb1_sq142 = xn2 & multm_reduce_sc142;
  assign multm_reduce_mulb1_sq143 = xn2 & multm_reduce_sc143;
  assign multm_reduce_mulb1_sq144 = xn2 & multm_reduce_sc144;
  assign multm_reduce_mulb1_sq145 = xn2 & multm_reduce_sc145;
  assign multm_reduce_mulb1_sq146 = xn2 & multm_reduce_sc146;
  assign multm_reduce_mulb1_sq147 = xn2 & multm_reduce_sc147;
  assign multm_reduce_mulb1_sq148 = xn2 & multm_reduce_sc148;
  assign multm_reduce_mulb1_sq149 = xn2 & multm_reduce_sc149;
  assign multm_reduce_mulb1_sq150 = xn2 & multm_reduce_sc150;
  assign multm_reduce_mulb1_sq151 = xn2 & multm_reduce_sc151;
  assign multm_reduce_mulb1_sq152 = xn2 & multm_reduce_sc152;
  assign multm_reduce_mulb1_sq153 = xn2 & multm_reduce_sc153;
  assign multm_reduce_mulb1_sq154 = xn2 & multm_reduce_sc154;
  assign multm_reduce_mulb1_sq155 = xn2 & multm_reduce_sc155;
  assign multm_reduce_mulb1_sq156 = xn2 & multm_reduce_sc156;
  assign multm_reduce_mulb1_sq157 = xn2 & multm_reduce_sc157;
  assign multm_reduce_mulb1_sq158 = xn2 & multm_reduce_sc158;
  assign multm_reduce_mulb1_sq159 = xn2 & multm_reduce_sc159;
  assign multm_reduce_mulb1_sq160 = xn2 & multm_reduce_sc160;
  assign multm_reduce_mulb1_sq161 = xn2 & multm_reduce_sc161;
  assign multm_reduce_mulb1_sq162 = xn2 & multm_reduce_sc162;
  assign multm_reduce_mulb1_sq163 = xn2 & multm_reduce_sc163;
  assign multm_reduce_mulb1_sq164 = xn2 & multm_reduce_sc164;
  assign multm_reduce_mulb1_sq165 = xn2 & multm_reduce_sc165;
  assign multm_reduce_mulb1_sq166 = xn2 & multm_reduce_sc166;
  assign multm_reduce_mulb1_sq167 = xn2 & multm_reduce_sc167;
  assign multm_reduce_mulb1_sq168 = xn2 & multm_reduce_sc168;
  assign multm_reduce_mulb1_sq169 = xn2 & multm_reduce_sc169;
  assign multm_reduce_mulb1_sq170 = xn2 & multm_reduce_sc170;
  assign multm_reduce_mulb1_sq171 = xn2 & multm_reduce_sc171;
  assign multm_reduce_mulb1_sq172 = xn2 & multm_reduce_sc172;
  assign multm_reduce_mulb1_sq173 = xn2 & multm_reduce_sc173;
  assign multm_reduce_mulb1_sq174 = xn2 & multm_reduce_sc174;
  assign multm_reduce_mulb1_sq175 = xn2 & multm_reduce_sc175;
  assign multm_reduce_mulb1_sq176 = xn2 & multm_reduce_sc176;
  assign multm_reduce_mulb1_sq177 = xn2 & multm_reduce_sc177;
  assign multm_reduce_mulb1_sq178 = xn2 & multm_reduce_sc178;
  assign multm_reduce_mulb1_sq179 = xn2 & multm_reduce_sc179;
  assign multm_reduce_mulb1_sq180 = xn2 & multm_reduce_sc180;
  assign multm_reduce_mulb1_sq181 = xn2 & multm_reduce_sc181;
  assign multm_reduce_mulb1_sq182 = xn2 & multm_reduce_sc182;
  assign multm_reduce_mulsc_mulb_add3_maj3_or3_wx = multm_reduce_mulsc_mulb_add3_maj3_wx | multm_reduce_mulsc_mulb_add3_maj3_wy;
  assign multm_reduce_mulsc_mulb_add3_maj3_wx = multm_reduce_mulsc_mulb_yoc183 & multm_reduce_mulsc_mulb_cq183;
  assign multm_reduce_mulsc_mulb_add3_maj3_wy = multm_reduce_mulsc_mulb_yoc183 & multm_reduce_mulsc_mulb_pc183;
  assign multm_reduce_mulsc_mulb_add3_maj3_xy = multm_reduce_mulsc_mulb_cq183 & multm_reduce_mulsc_mulb_pc183;
  assign multm_reduce_mulsc_mulb_add3_xor3_wx = multm_reduce_mulsc_mulb_yoc183 ^ multm_reduce_mulsc_mulb_cq183;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx0 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx0 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy0;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx1 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx1 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy1;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx2 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx2 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy2;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx3 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx3 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy3;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx4 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx4 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy4;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx5 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx5 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy5;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx6 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx6 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy6;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx7 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx7 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy7;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx8 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx8 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy8;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx9 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx9 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy9;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx10 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx10 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy10;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx11 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx11 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy11;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx12 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx12 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy12;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx13 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx13 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy13;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx14 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx14 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy14;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx15 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx15 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy15;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx16 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx16 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy16;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx17 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx17 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy17;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx18 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx18 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy18;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx19 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx19 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy19;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx20 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx20 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy20;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx21 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx21 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy21;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx22 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx22 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy22;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx23 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx23 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy23;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx24 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx24 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy24;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx25 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx25 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy25;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx26 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx26 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy26;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx27 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx27 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy27;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx28 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx28 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy28;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx29 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx29 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy29;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx30 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx30 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy30;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx31 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx31 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy31;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx32 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx32 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy32;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx33 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx33 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy33;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx34 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx34 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy34;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx35 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx35 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy35;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx36 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx36 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy36;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx37 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx37 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy37;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx38 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx38 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy38;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx39 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx39 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy39;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx40 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx40 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy40;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx41 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx41 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy41;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx42 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx42 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy42;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx43 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx43 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy43;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx44 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx44 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy44;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx45 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx45 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy45;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx46 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx46 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy46;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx47 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx47 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy47;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx48 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx48 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy48;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx49 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx49 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy49;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx50 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx50 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy50;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx51 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx51 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy51;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx52 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx52 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy52;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx53 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx53 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy53;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx54 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx54 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy54;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx55 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx55 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy55;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx56 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx56 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy56;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx57 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx57 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy57;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx58 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx58 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy58;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx59 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx59 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy59;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx60 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx60 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy60;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx61 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx61 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy61;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx62 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx62 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy62;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx63 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx63 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy63;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx64 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx64 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy64;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx65 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx65 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy65;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx66 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx66 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy66;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx67 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx67 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy67;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx68 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx68 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy68;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx69 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx69 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy69;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx70 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx70 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy70;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx71 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx71 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy71;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx72 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx72 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy72;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx73 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx73 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy73;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx74 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx74 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy74;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx75 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx75 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy75;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx76 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx76 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy76;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx77 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx77 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy77;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx78 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx78 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy78;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx79 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx79 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy79;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx80 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx80 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy80;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx81 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx81 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy81;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx82 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx82 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy82;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx83 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx83 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy83;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx84 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx84 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy84;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx85 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx85 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy85;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx86 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx86 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy86;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx87 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx87 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy87;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx88 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx88 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy88;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx89 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx89 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy89;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx90 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx90 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy90;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx91 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx91 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy91;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx92 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx92 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy92;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx93 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx93 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy93;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx94 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx94 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy94;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx95 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx95 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy95;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx96 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx96 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy96;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx97 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx97 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy97;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx98 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx98 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy98;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx99 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx99 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy99;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx100 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx100 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy100;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx101 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx101 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy101;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx102 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx102 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy102;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx103 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx103 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy103;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx104 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx104 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy104;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx105 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx105 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy105;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx106 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx106 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy106;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx107 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx107 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy107;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx108 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx108 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy108;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx109 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx109 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy109;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx110 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx110 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy110;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx111 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx111 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy111;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx112 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx112 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy112;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx113 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx113 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy113;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx114 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx114 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy114;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx115 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx115 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy115;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx116 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx116 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy116;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx117 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx117 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy117;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx118 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx118 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy118;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx119 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx119 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy119;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx120 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx120 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy120;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx121 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx121 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy121;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx122 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx122 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy122;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx123 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx123 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy123;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx124 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx124 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy124;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx125 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx125 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy125;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx126 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx126 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy126;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx127 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx127 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy127;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx128 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx128 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy128;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx129 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx129 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy129;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx130 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx130 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy130;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx131 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx131 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy131;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx132 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx132 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy132;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx133 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx133 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy133;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx134 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx134 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy134;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx135 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx135 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy135;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx136 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx136 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy136;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx137 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx137 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy137;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx138 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx138 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy138;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx139 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx139 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy139;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx140 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx140 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy140;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx141 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx141 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy141;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx142 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx142 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy142;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx143 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx143 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy143;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx144 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx144 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy144;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx145 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx145 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy145;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx146 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx146 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy146;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx147 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx147 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy147;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx148 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx148 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy148;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx149 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx149 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy149;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx150 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx150 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy150;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx151 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx151 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy151;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx152 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx152 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy152;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx153 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx153 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy153;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx154 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx154 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy154;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx155 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx155 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy155;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx156 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx156 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy156;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx157 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx157 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy157;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx158 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx158 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy158;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx159 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx159 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy159;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx160 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx160 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy160;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx161 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx161 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy161;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx162 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx162 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy162;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx163 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx163 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy163;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx164 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx164 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy164;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx165 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx165 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy165;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx166 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx166 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy166;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx167 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx167 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy167;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx168 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx168 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy168;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx169 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx169 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy169;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx170 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx170 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy170;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx171 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx171 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy171;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx172 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx172 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy172;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx173 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx173 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy173;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx174 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx174 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy174;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx175 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx175 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy175;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx176 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx176 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy176;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx177 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx177 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy177;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx178 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx178 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy178;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx179 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx179 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy179;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx180 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx180 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy180;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx181 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx181 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy181;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx182 = multm_reduce_mulsc_mulb_add3b0_maj3b_wx182 | multm_reduce_mulsc_mulb_add3b0_maj3b_wy182;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx0 = multm_reduce_mulsc_mulb_sq1 & multm_reduce_mulsc_mulb_cq0;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx1 = multm_reduce_mulsc_mulb_sq2 & multm_reduce_mulsc_mulb_cq1;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx2 = multm_reduce_mulsc_mulb_sq3 & multm_reduce_mulsc_mulb_cq2;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx3 = multm_reduce_mulsc_mulb_sq4 & multm_reduce_mulsc_mulb_cq3;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx4 = multm_reduce_mulsc_mulb_sq5 & multm_reduce_mulsc_mulb_cq4;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx5 = multm_reduce_mulsc_mulb_sq6 & multm_reduce_mulsc_mulb_cq5;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx6 = multm_reduce_mulsc_mulb_sq7 & multm_reduce_mulsc_mulb_cq6;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx7 = multm_reduce_mulsc_mulb_sq8 & multm_reduce_mulsc_mulb_cq7;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx8 = multm_reduce_mulsc_mulb_sq9 & multm_reduce_mulsc_mulb_cq8;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx9 = multm_reduce_mulsc_mulb_sq10 & multm_reduce_mulsc_mulb_cq9;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx10 = multm_reduce_mulsc_mulb_sq11 & multm_reduce_mulsc_mulb_cq10;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx11 = multm_reduce_mulsc_mulb_sq12 & multm_reduce_mulsc_mulb_cq11;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx12 = multm_reduce_mulsc_mulb_sq13 & multm_reduce_mulsc_mulb_cq12;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx13 = multm_reduce_mulsc_mulb_sq14 & multm_reduce_mulsc_mulb_cq13;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx14 = multm_reduce_mulsc_mulb_sq15 & multm_reduce_mulsc_mulb_cq14;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx15 = multm_reduce_mulsc_mulb_sq16 & multm_reduce_mulsc_mulb_cq15;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx16 = multm_reduce_mulsc_mulb_sq17 & multm_reduce_mulsc_mulb_cq16;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx17 = multm_reduce_mulsc_mulb_sq18 & multm_reduce_mulsc_mulb_cq17;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx18 = multm_reduce_mulsc_mulb_sq19 & multm_reduce_mulsc_mulb_cq18;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx19 = multm_reduce_mulsc_mulb_sq20 & multm_reduce_mulsc_mulb_cq19;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx20 = multm_reduce_mulsc_mulb_sq21 & multm_reduce_mulsc_mulb_cq20;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx21 = multm_reduce_mulsc_mulb_sq22 & multm_reduce_mulsc_mulb_cq21;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx22 = multm_reduce_mulsc_mulb_sq23 & multm_reduce_mulsc_mulb_cq22;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx23 = multm_reduce_mulsc_mulb_sq24 & multm_reduce_mulsc_mulb_cq23;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx24 = multm_reduce_mulsc_mulb_sq25 & multm_reduce_mulsc_mulb_cq24;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx25 = multm_reduce_mulsc_mulb_sq26 & multm_reduce_mulsc_mulb_cq25;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx26 = multm_reduce_mulsc_mulb_sq27 & multm_reduce_mulsc_mulb_cq26;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx27 = multm_reduce_mulsc_mulb_sq28 & multm_reduce_mulsc_mulb_cq27;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx28 = multm_reduce_mulsc_mulb_sq29 & multm_reduce_mulsc_mulb_cq28;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx29 = multm_reduce_mulsc_mulb_sq30 & multm_reduce_mulsc_mulb_cq29;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx30 = multm_reduce_mulsc_mulb_sq31 & multm_reduce_mulsc_mulb_cq30;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx31 = multm_reduce_mulsc_mulb_sq32 & multm_reduce_mulsc_mulb_cq31;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx32 = multm_reduce_mulsc_mulb_sq33 & multm_reduce_mulsc_mulb_cq32;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx33 = multm_reduce_mulsc_mulb_sq34 & multm_reduce_mulsc_mulb_cq33;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx34 = multm_reduce_mulsc_mulb_sq35 & multm_reduce_mulsc_mulb_cq34;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx35 = multm_reduce_mulsc_mulb_sq36 & multm_reduce_mulsc_mulb_cq35;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx36 = multm_reduce_mulsc_mulb_sq37 & multm_reduce_mulsc_mulb_cq36;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx37 = multm_reduce_mulsc_mulb_sq38 & multm_reduce_mulsc_mulb_cq37;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx38 = multm_reduce_mulsc_mulb_sq39 & multm_reduce_mulsc_mulb_cq38;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx39 = multm_reduce_mulsc_mulb_sq40 & multm_reduce_mulsc_mulb_cq39;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx40 = multm_reduce_mulsc_mulb_sq41 & multm_reduce_mulsc_mulb_cq40;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx41 = multm_reduce_mulsc_mulb_sq42 & multm_reduce_mulsc_mulb_cq41;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx42 = multm_reduce_mulsc_mulb_sq43 & multm_reduce_mulsc_mulb_cq42;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx43 = multm_reduce_mulsc_mulb_sq44 & multm_reduce_mulsc_mulb_cq43;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx44 = multm_reduce_mulsc_mulb_sq45 & multm_reduce_mulsc_mulb_cq44;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx45 = multm_reduce_mulsc_mulb_sq46 & multm_reduce_mulsc_mulb_cq45;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx46 = multm_reduce_mulsc_mulb_sq47 & multm_reduce_mulsc_mulb_cq46;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx47 = multm_reduce_mulsc_mulb_sq48 & multm_reduce_mulsc_mulb_cq47;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx48 = multm_reduce_mulsc_mulb_sq49 & multm_reduce_mulsc_mulb_cq48;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx49 = multm_reduce_mulsc_mulb_sq50 & multm_reduce_mulsc_mulb_cq49;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx50 = multm_reduce_mulsc_mulb_sq51 & multm_reduce_mulsc_mulb_cq50;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx51 = multm_reduce_mulsc_mulb_sq52 & multm_reduce_mulsc_mulb_cq51;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx52 = multm_reduce_mulsc_mulb_sq53 & multm_reduce_mulsc_mulb_cq52;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx53 = multm_reduce_mulsc_mulb_sq54 & multm_reduce_mulsc_mulb_cq53;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx54 = multm_reduce_mulsc_mulb_sq55 & multm_reduce_mulsc_mulb_cq54;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx55 = multm_reduce_mulsc_mulb_sq56 & multm_reduce_mulsc_mulb_cq55;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx56 = multm_reduce_mulsc_mulb_sq57 & multm_reduce_mulsc_mulb_cq56;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx57 = multm_reduce_mulsc_mulb_sq58 & multm_reduce_mulsc_mulb_cq57;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx58 = multm_reduce_mulsc_mulb_sq59 & multm_reduce_mulsc_mulb_cq58;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx59 = multm_reduce_mulsc_mulb_sq60 & multm_reduce_mulsc_mulb_cq59;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx60 = multm_reduce_mulsc_mulb_sq61 & multm_reduce_mulsc_mulb_cq60;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx61 = multm_reduce_mulsc_mulb_sq62 & multm_reduce_mulsc_mulb_cq61;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx62 = multm_reduce_mulsc_mulb_sq63 & multm_reduce_mulsc_mulb_cq62;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx63 = multm_reduce_mulsc_mulb_sq64 & multm_reduce_mulsc_mulb_cq63;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx64 = multm_reduce_mulsc_mulb_sq65 & multm_reduce_mulsc_mulb_cq64;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx65 = multm_reduce_mulsc_mulb_sq66 & multm_reduce_mulsc_mulb_cq65;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx66 = multm_reduce_mulsc_mulb_sq67 & multm_reduce_mulsc_mulb_cq66;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx67 = multm_reduce_mulsc_mulb_sq68 & multm_reduce_mulsc_mulb_cq67;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx68 = multm_reduce_mulsc_mulb_sq69 & multm_reduce_mulsc_mulb_cq68;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx69 = multm_reduce_mulsc_mulb_sq70 & multm_reduce_mulsc_mulb_cq69;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx70 = multm_reduce_mulsc_mulb_sq71 & multm_reduce_mulsc_mulb_cq70;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx71 = multm_reduce_mulsc_mulb_sq72 & multm_reduce_mulsc_mulb_cq71;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx72 = multm_reduce_mulsc_mulb_sq73 & multm_reduce_mulsc_mulb_cq72;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx73 = multm_reduce_mulsc_mulb_sq74 & multm_reduce_mulsc_mulb_cq73;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx74 = multm_reduce_mulsc_mulb_sq75 & multm_reduce_mulsc_mulb_cq74;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx75 = multm_reduce_mulsc_mulb_sq76 & multm_reduce_mulsc_mulb_cq75;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx76 = multm_reduce_mulsc_mulb_sq77 & multm_reduce_mulsc_mulb_cq76;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx77 = multm_reduce_mulsc_mulb_sq78 & multm_reduce_mulsc_mulb_cq77;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx78 = multm_reduce_mulsc_mulb_sq79 & multm_reduce_mulsc_mulb_cq78;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx79 = multm_reduce_mulsc_mulb_sq80 & multm_reduce_mulsc_mulb_cq79;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx80 = multm_reduce_mulsc_mulb_sq81 & multm_reduce_mulsc_mulb_cq80;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx81 = multm_reduce_mulsc_mulb_sq82 & multm_reduce_mulsc_mulb_cq81;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx82 = multm_reduce_mulsc_mulb_sq83 & multm_reduce_mulsc_mulb_cq82;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx83 = multm_reduce_mulsc_mulb_sq84 & multm_reduce_mulsc_mulb_cq83;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx84 = multm_reduce_mulsc_mulb_sq85 & multm_reduce_mulsc_mulb_cq84;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx85 = multm_reduce_mulsc_mulb_sq86 & multm_reduce_mulsc_mulb_cq85;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx86 = multm_reduce_mulsc_mulb_sq87 & multm_reduce_mulsc_mulb_cq86;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx87 = multm_reduce_mulsc_mulb_sq88 & multm_reduce_mulsc_mulb_cq87;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx88 = multm_reduce_mulsc_mulb_sq89 & multm_reduce_mulsc_mulb_cq88;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx89 = multm_reduce_mulsc_mulb_sq90 & multm_reduce_mulsc_mulb_cq89;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx90 = multm_reduce_mulsc_mulb_sq91 & multm_reduce_mulsc_mulb_cq90;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx91 = multm_reduce_mulsc_mulb_sq92 & multm_reduce_mulsc_mulb_cq91;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx92 = multm_reduce_mulsc_mulb_sq93 & multm_reduce_mulsc_mulb_cq92;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx93 = multm_reduce_mulsc_mulb_sq94 & multm_reduce_mulsc_mulb_cq93;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx94 = multm_reduce_mulsc_mulb_sq95 & multm_reduce_mulsc_mulb_cq94;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx95 = multm_reduce_mulsc_mulb_sq96 & multm_reduce_mulsc_mulb_cq95;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx96 = multm_reduce_mulsc_mulb_sq97 & multm_reduce_mulsc_mulb_cq96;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx97 = multm_reduce_mulsc_mulb_sq98 & multm_reduce_mulsc_mulb_cq97;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx98 = multm_reduce_mulsc_mulb_sq99 & multm_reduce_mulsc_mulb_cq98;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx99 = multm_reduce_mulsc_mulb_sq100 & multm_reduce_mulsc_mulb_cq99;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx100 = multm_reduce_mulsc_mulb_sq101 & multm_reduce_mulsc_mulb_cq100;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx101 = multm_reduce_mulsc_mulb_sq102 & multm_reduce_mulsc_mulb_cq101;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx102 = multm_reduce_mulsc_mulb_sq103 & multm_reduce_mulsc_mulb_cq102;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx103 = multm_reduce_mulsc_mulb_sq104 & multm_reduce_mulsc_mulb_cq103;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx104 = multm_reduce_mulsc_mulb_sq105 & multm_reduce_mulsc_mulb_cq104;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx105 = multm_reduce_mulsc_mulb_sq106 & multm_reduce_mulsc_mulb_cq105;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx106 = multm_reduce_mulsc_mulb_sq107 & multm_reduce_mulsc_mulb_cq106;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx107 = multm_reduce_mulsc_mulb_sq108 & multm_reduce_mulsc_mulb_cq107;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx108 = multm_reduce_mulsc_mulb_sq109 & multm_reduce_mulsc_mulb_cq108;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx109 = multm_reduce_mulsc_mulb_sq110 & multm_reduce_mulsc_mulb_cq109;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx110 = multm_reduce_mulsc_mulb_sq111 & multm_reduce_mulsc_mulb_cq110;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx111 = multm_reduce_mulsc_mulb_sq112 & multm_reduce_mulsc_mulb_cq111;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx112 = multm_reduce_mulsc_mulb_sq113 & multm_reduce_mulsc_mulb_cq112;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx113 = multm_reduce_mulsc_mulb_sq114 & multm_reduce_mulsc_mulb_cq113;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx114 = multm_reduce_mulsc_mulb_sq115 & multm_reduce_mulsc_mulb_cq114;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx115 = multm_reduce_mulsc_mulb_sq116 & multm_reduce_mulsc_mulb_cq115;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx116 = multm_reduce_mulsc_mulb_sq117 & multm_reduce_mulsc_mulb_cq116;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx117 = multm_reduce_mulsc_mulb_sq118 & multm_reduce_mulsc_mulb_cq117;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx118 = multm_reduce_mulsc_mulb_sq119 & multm_reduce_mulsc_mulb_cq118;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx119 = multm_reduce_mulsc_mulb_sq120 & multm_reduce_mulsc_mulb_cq119;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx120 = multm_reduce_mulsc_mulb_sq121 & multm_reduce_mulsc_mulb_cq120;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx121 = multm_reduce_mulsc_mulb_sq122 & multm_reduce_mulsc_mulb_cq121;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx122 = multm_reduce_mulsc_mulb_sq123 & multm_reduce_mulsc_mulb_cq122;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx123 = multm_reduce_mulsc_mulb_sq124 & multm_reduce_mulsc_mulb_cq123;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx124 = multm_reduce_mulsc_mulb_sq125 & multm_reduce_mulsc_mulb_cq124;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx125 = multm_reduce_mulsc_mulb_sq126 & multm_reduce_mulsc_mulb_cq125;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx126 = multm_reduce_mulsc_mulb_sq127 & multm_reduce_mulsc_mulb_cq126;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx127 = multm_reduce_mulsc_mulb_sq128 & multm_reduce_mulsc_mulb_cq127;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx128 = multm_reduce_mulsc_mulb_sq129 & multm_reduce_mulsc_mulb_cq128;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx129 = multm_reduce_mulsc_mulb_sq130 & multm_reduce_mulsc_mulb_cq129;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx130 = multm_reduce_mulsc_mulb_sq131 & multm_reduce_mulsc_mulb_cq130;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx131 = multm_reduce_mulsc_mulb_sq132 & multm_reduce_mulsc_mulb_cq131;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx132 = multm_reduce_mulsc_mulb_sq133 & multm_reduce_mulsc_mulb_cq132;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx133 = multm_reduce_mulsc_mulb_sq134 & multm_reduce_mulsc_mulb_cq133;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx134 = multm_reduce_mulsc_mulb_sq135 & multm_reduce_mulsc_mulb_cq134;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx135 = multm_reduce_mulsc_mulb_sq136 & multm_reduce_mulsc_mulb_cq135;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx136 = multm_reduce_mulsc_mulb_sq137 & multm_reduce_mulsc_mulb_cq136;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx137 = multm_reduce_mulsc_mulb_sq138 & multm_reduce_mulsc_mulb_cq137;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx138 = multm_reduce_mulsc_mulb_sq139 & multm_reduce_mulsc_mulb_cq138;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx139 = multm_reduce_mulsc_mulb_sq140 & multm_reduce_mulsc_mulb_cq139;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx140 = multm_reduce_mulsc_mulb_sq141 & multm_reduce_mulsc_mulb_cq140;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx141 = multm_reduce_mulsc_mulb_sq142 & multm_reduce_mulsc_mulb_cq141;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx142 = multm_reduce_mulsc_mulb_sq143 & multm_reduce_mulsc_mulb_cq142;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx143 = multm_reduce_mulsc_mulb_sq144 & multm_reduce_mulsc_mulb_cq143;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx144 = multm_reduce_mulsc_mulb_sq145 & multm_reduce_mulsc_mulb_cq144;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx145 = multm_reduce_mulsc_mulb_sq146 & multm_reduce_mulsc_mulb_cq145;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx146 = multm_reduce_mulsc_mulb_sq147 & multm_reduce_mulsc_mulb_cq146;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx147 = multm_reduce_mulsc_mulb_sq148 & multm_reduce_mulsc_mulb_cq147;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx148 = multm_reduce_mulsc_mulb_sq149 & multm_reduce_mulsc_mulb_cq148;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx149 = multm_reduce_mulsc_mulb_sq150 & multm_reduce_mulsc_mulb_cq149;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx150 = multm_reduce_mulsc_mulb_sq151 & multm_reduce_mulsc_mulb_cq150;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx151 = multm_reduce_mulsc_mulb_sq152 & multm_reduce_mulsc_mulb_cq151;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx152 = multm_reduce_mulsc_mulb_sq153 & multm_reduce_mulsc_mulb_cq152;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx153 = multm_reduce_mulsc_mulb_sq154 & multm_reduce_mulsc_mulb_cq153;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx154 = multm_reduce_mulsc_mulb_sq155 & multm_reduce_mulsc_mulb_cq154;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx155 = multm_reduce_mulsc_mulb_sq156 & multm_reduce_mulsc_mulb_cq155;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx156 = multm_reduce_mulsc_mulb_sq157 & multm_reduce_mulsc_mulb_cq156;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx157 = multm_reduce_mulsc_mulb_sq158 & multm_reduce_mulsc_mulb_cq157;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx158 = multm_reduce_mulsc_mulb_sq159 & multm_reduce_mulsc_mulb_cq158;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx159 = multm_reduce_mulsc_mulb_sq160 & multm_reduce_mulsc_mulb_cq159;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx160 = multm_reduce_mulsc_mulb_sq161 & multm_reduce_mulsc_mulb_cq160;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx161 = multm_reduce_mulsc_mulb_sq162 & multm_reduce_mulsc_mulb_cq161;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx162 = multm_reduce_mulsc_mulb_sq163 & multm_reduce_mulsc_mulb_cq162;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx163 = multm_reduce_mulsc_mulb_sq164 & multm_reduce_mulsc_mulb_cq163;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx164 = multm_reduce_mulsc_mulb_sq165 & multm_reduce_mulsc_mulb_cq164;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx165 = multm_reduce_mulsc_mulb_sq166 & multm_reduce_mulsc_mulb_cq165;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx166 = multm_reduce_mulsc_mulb_sq167 & multm_reduce_mulsc_mulb_cq166;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx167 = multm_reduce_mulsc_mulb_sq168 & multm_reduce_mulsc_mulb_cq167;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx168 = multm_reduce_mulsc_mulb_sq169 & multm_reduce_mulsc_mulb_cq168;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx169 = multm_reduce_mulsc_mulb_sq170 & multm_reduce_mulsc_mulb_cq169;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx170 = multm_reduce_mulsc_mulb_sq171 & multm_reduce_mulsc_mulb_cq170;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx171 = multm_reduce_mulsc_mulb_sq172 & multm_reduce_mulsc_mulb_cq171;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx172 = multm_reduce_mulsc_mulb_sq173 & multm_reduce_mulsc_mulb_cq172;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx173 = multm_reduce_mulsc_mulb_sq174 & multm_reduce_mulsc_mulb_cq173;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx174 = multm_reduce_mulsc_mulb_sq175 & multm_reduce_mulsc_mulb_cq174;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx175 = multm_reduce_mulsc_mulb_sq176 & multm_reduce_mulsc_mulb_cq175;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx176 = multm_reduce_mulsc_mulb_sq177 & multm_reduce_mulsc_mulb_cq176;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx177 = multm_reduce_mulsc_mulb_sq178 & multm_reduce_mulsc_mulb_cq177;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx178 = multm_reduce_mulsc_mulb_sq179 & multm_reduce_mulsc_mulb_cq178;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx179 = multm_reduce_mulsc_mulb_sq180 & multm_reduce_mulsc_mulb_cq179;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx180 = multm_reduce_mulsc_mulb_sq181 & multm_reduce_mulsc_mulb_cq180;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx181 = multm_reduce_mulsc_mulb_sq182 & multm_reduce_mulsc_mulb_cq181;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wx182 = multm_reduce_mulsc_mulb_sq183 & multm_reduce_mulsc_mulb_cq182;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy0 = multm_reduce_mulsc_mulb_sq1 & multm_reduce_mulsc_mulb_yos1;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy1 = multm_reduce_mulsc_mulb_sq2 & multm_reduce_mulsc_mulb_yos2;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy2 = multm_reduce_mulsc_mulb_sq3 & multm_reduce_mulsc_mulb_yos3;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy3 = multm_reduce_mulsc_mulb_sq4 & multm_reduce_mulsc_mulb_yos4;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy4 = multm_reduce_mulsc_mulb_sq5 & multm_reduce_mulsc_mulb_yos5;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy5 = multm_reduce_mulsc_mulb_sq6 & multm_reduce_mulsc_mulb_yos6;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy6 = multm_reduce_mulsc_mulb_sq7 & multm_reduce_mulsc_mulb_yos7;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy7 = multm_reduce_mulsc_mulb_sq8 & multm_reduce_mulsc_mulb_yos8;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy8 = multm_reduce_mulsc_mulb_sq9 & multm_reduce_mulsc_mulb_yos9;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy9 = multm_reduce_mulsc_mulb_sq10 & multm_reduce_mulsc_mulb_yos10;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy10 = multm_reduce_mulsc_mulb_sq11 & multm_reduce_mulsc_mulb_yos11;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy11 = multm_reduce_mulsc_mulb_sq12 & multm_reduce_mulsc_mulb_yos12;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy12 = multm_reduce_mulsc_mulb_sq13 & multm_reduce_mulsc_mulb_yos13;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy13 = multm_reduce_mulsc_mulb_sq14 & multm_reduce_mulsc_mulb_yos14;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy14 = multm_reduce_mulsc_mulb_sq15 & multm_reduce_mulsc_mulb_yos15;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy15 = multm_reduce_mulsc_mulb_sq16 & multm_reduce_mulsc_mulb_yos16;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy16 = multm_reduce_mulsc_mulb_sq17 & multm_reduce_mulsc_mulb_yos17;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy17 = multm_reduce_mulsc_mulb_sq18 & multm_reduce_mulsc_mulb_yos18;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy18 = multm_reduce_mulsc_mulb_sq19 & multm_reduce_mulsc_mulb_yos19;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy19 = multm_reduce_mulsc_mulb_sq20 & multm_reduce_mulsc_mulb_yos20;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy20 = multm_reduce_mulsc_mulb_sq21 & multm_reduce_mulsc_mulb_yos21;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy21 = multm_reduce_mulsc_mulb_sq22 & multm_reduce_mulsc_mulb_yos22;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy22 = multm_reduce_mulsc_mulb_sq23 & multm_reduce_mulsc_mulb_yos23;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy23 = multm_reduce_mulsc_mulb_sq24 & multm_reduce_mulsc_mulb_yos24;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy24 = multm_reduce_mulsc_mulb_sq25 & multm_reduce_mulsc_mulb_yos25;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy25 = multm_reduce_mulsc_mulb_sq26 & multm_reduce_mulsc_mulb_yos26;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy26 = multm_reduce_mulsc_mulb_sq27 & multm_reduce_mulsc_mulb_yos27;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy27 = multm_reduce_mulsc_mulb_sq28 & multm_reduce_mulsc_mulb_yos28;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy28 = multm_reduce_mulsc_mulb_sq29 & multm_reduce_mulsc_mulb_yos29;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy29 = multm_reduce_mulsc_mulb_sq30 & multm_reduce_mulsc_mulb_yos30;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy30 = multm_reduce_mulsc_mulb_sq31 & multm_reduce_mulsc_mulb_yos31;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy31 = multm_reduce_mulsc_mulb_sq32 & multm_reduce_mulsc_mulb_yos32;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy32 = multm_reduce_mulsc_mulb_sq33 & multm_reduce_mulsc_mulb_yos33;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy33 = multm_reduce_mulsc_mulb_sq34 & multm_reduce_mulsc_mulb_yos34;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy34 = multm_reduce_mulsc_mulb_sq35 & multm_reduce_mulsc_mulb_yos35;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy35 = multm_reduce_mulsc_mulb_sq36 & multm_reduce_mulsc_mulb_yos36;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy36 = multm_reduce_mulsc_mulb_sq37 & multm_reduce_mulsc_mulb_yos37;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy37 = multm_reduce_mulsc_mulb_sq38 & multm_reduce_mulsc_mulb_yos38;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy38 = multm_reduce_mulsc_mulb_sq39 & multm_reduce_mulsc_mulb_yos39;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy39 = multm_reduce_mulsc_mulb_sq40 & multm_reduce_mulsc_mulb_yos40;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy40 = multm_reduce_mulsc_mulb_sq41 & multm_reduce_mulsc_mulb_yos41;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy41 = multm_reduce_mulsc_mulb_sq42 & multm_reduce_mulsc_mulb_yos42;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy42 = multm_reduce_mulsc_mulb_sq43 & multm_reduce_mulsc_mulb_yos43;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy43 = multm_reduce_mulsc_mulb_sq44 & multm_reduce_mulsc_mulb_yos44;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy44 = multm_reduce_mulsc_mulb_sq45 & multm_reduce_mulsc_mulb_yos45;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy45 = multm_reduce_mulsc_mulb_sq46 & multm_reduce_mulsc_mulb_yos46;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy46 = multm_reduce_mulsc_mulb_sq47 & multm_reduce_mulsc_mulb_yos47;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy47 = multm_reduce_mulsc_mulb_sq48 & multm_reduce_mulsc_mulb_yos48;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy48 = multm_reduce_mulsc_mulb_sq49 & multm_reduce_mulsc_mulb_yos49;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy49 = multm_reduce_mulsc_mulb_sq50 & multm_reduce_mulsc_mulb_yos50;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy50 = multm_reduce_mulsc_mulb_sq51 & multm_reduce_mulsc_mulb_yos51;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy51 = multm_reduce_mulsc_mulb_sq52 & multm_reduce_mulsc_mulb_yos52;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy52 = multm_reduce_mulsc_mulb_sq53 & multm_reduce_mulsc_mulb_yos53;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy53 = multm_reduce_mulsc_mulb_sq54 & multm_reduce_mulsc_mulb_yos54;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy54 = multm_reduce_mulsc_mulb_sq55 & multm_reduce_mulsc_mulb_yos55;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy55 = multm_reduce_mulsc_mulb_sq56 & multm_reduce_mulsc_mulb_yos56;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy56 = multm_reduce_mulsc_mulb_sq57 & multm_reduce_mulsc_mulb_yos57;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy57 = multm_reduce_mulsc_mulb_sq58 & multm_reduce_mulsc_mulb_yos58;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy58 = multm_reduce_mulsc_mulb_sq59 & multm_reduce_mulsc_mulb_yos59;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy59 = multm_reduce_mulsc_mulb_sq60 & multm_reduce_mulsc_mulb_yos60;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy60 = multm_reduce_mulsc_mulb_sq61 & multm_reduce_mulsc_mulb_yos61;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy61 = multm_reduce_mulsc_mulb_sq62 & multm_reduce_mulsc_mulb_yos62;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy62 = multm_reduce_mulsc_mulb_sq63 & multm_reduce_mulsc_mulb_yos63;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy63 = multm_reduce_mulsc_mulb_sq64 & multm_reduce_mulsc_mulb_yos64;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy64 = multm_reduce_mulsc_mulb_sq65 & multm_reduce_mulsc_mulb_yos65;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy65 = multm_reduce_mulsc_mulb_sq66 & multm_reduce_mulsc_mulb_yos66;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy66 = multm_reduce_mulsc_mulb_sq67 & multm_reduce_mulsc_mulb_yos67;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy67 = multm_reduce_mulsc_mulb_sq68 & multm_reduce_mulsc_mulb_yos68;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy68 = multm_reduce_mulsc_mulb_sq69 & multm_reduce_mulsc_mulb_yos69;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy69 = multm_reduce_mulsc_mulb_sq70 & multm_reduce_mulsc_mulb_yos70;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy70 = multm_reduce_mulsc_mulb_sq71 & multm_reduce_mulsc_mulb_yos71;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy71 = multm_reduce_mulsc_mulb_sq72 & multm_reduce_mulsc_mulb_yos72;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy72 = multm_reduce_mulsc_mulb_sq73 & multm_reduce_mulsc_mulb_yos73;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy73 = multm_reduce_mulsc_mulb_sq74 & multm_reduce_mulsc_mulb_yos74;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy74 = multm_reduce_mulsc_mulb_sq75 & multm_reduce_mulsc_mulb_yos75;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy75 = multm_reduce_mulsc_mulb_sq76 & multm_reduce_mulsc_mulb_yos76;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy76 = multm_reduce_mulsc_mulb_sq77 & multm_reduce_mulsc_mulb_yos77;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy77 = multm_reduce_mulsc_mulb_sq78 & multm_reduce_mulsc_mulb_yos78;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy78 = multm_reduce_mulsc_mulb_sq79 & multm_reduce_mulsc_mulb_yos79;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy79 = multm_reduce_mulsc_mulb_sq80 & multm_reduce_mulsc_mulb_yos80;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy80 = multm_reduce_mulsc_mulb_sq81 & multm_reduce_mulsc_mulb_yos81;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy81 = multm_reduce_mulsc_mulb_sq82 & multm_reduce_mulsc_mulb_yos82;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy82 = multm_reduce_mulsc_mulb_sq83 & multm_reduce_mulsc_mulb_yos83;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy83 = multm_reduce_mulsc_mulb_sq84 & multm_reduce_mulsc_mulb_yos84;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy84 = multm_reduce_mulsc_mulb_sq85 & multm_reduce_mulsc_mulb_yos85;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy85 = multm_reduce_mulsc_mulb_sq86 & multm_reduce_mulsc_mulb_yos86;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy86 = multm_reduce_mulsc_mulb_sq87 & multm_reduce_mulsc_mulb_yos87;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy87 = multm_reduce_mulsc_mulb_sq88 & multm_reduce_mulsc_mulb_yos88;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy88 = multm_reduce_mulsc_mulb_sq89 & multm_reduce_mulsc_mulb_yos89;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy89 = multm_reduce_mulsc_mulb_sq90 & multm_reduce_mulsc_mulb_yos90;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy90 = multm_reduce_mulsc_mulb_sq91 & multm_reduce_mulsc_mulb_yos91;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy91 = multm_reduce_mulsc_mulb_sq92 & multm_reduce_mulsc_mulb_yos92;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy92 = multm_reduce_mulsc_mulb_sq93 & multm_reduce_mulsc_mulb_yos93;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy93 = multm_reduce_mulsc_mulb_sq94 & multm_reduce_mulsc_mulb_yos94;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy94 = multm_reduce_mulsc_mulb_sq95 & multm_reduce_mulsc_mulb_yos95;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy95 = multm_reduce_mulsc_mulb_sq96 & multm_reduce_mulsc_mulb_yos96;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy96 = multm_reduce_mulsc_mulb_sq97 & multm_reduce_mulsc_mulb_yos97;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy97 = multm_reduce_mulsc_mulb_sq98 & multm_reduce_mulsc_mulb_yos98;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy98 = multm_reduce_mulsc_mulb_sq99 & multm_reduce_mulsc_mulb_yos99;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy99 = multm_reduce_mulsc_mulb_sq100 & multm_reduce_mulsc_mulb_yos100;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy100 = multm_reduce_mulsc_mulb_sq101 & multm_reduce_mulsc_mulb_yos101;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy101 = multm_reduce_mulsc_mulb_sq102 & multm_reduce_mulsc_mulb_yos102;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy102 = multm_reduce_mulsc_mulb_sq103 & multm_reduce_mulsc_mulb_yos103;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy103 = multm_reduce_mulsc_mulb_sq104 & multm_reduce_mulsc_mulb_yos104;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy104 = multm_reduce_mulsc_mulb_sq105 & multm_reduce_mulsc_mulb_yos105;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy105 = multm_reduce_mulsc_mulb_sq106 & multm_reduce_mulsc_mulb_yos106;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy106 = multm_reduce_mulsc_mulb_sq107 & multm_reduce_mulsc_mulb_yos107;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy107 = multm_reduce_mulsc_mulb_sq108 & multm_reduce_mulsc_mulb_yos108;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy108 = multm_reduce_mulsc_mulb_sq109 & multm_reduce_mulsc_mulb_yos109;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy109 = multm_reduce_mulsc_mulb_sq110 & multm_reduce_mulsc_mulb_yos110;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy110 = multm_reduce_mulsc_mulb_sq111 & multm_reduce_mulsc_mulb_yos111;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy111 = multm_reduce_mulsc_mulb_sq112 & multm_reduce_mulsc_mulb_yos112;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy112 = multm_reduce_mulsc_mulb_sq113 & multm_reduce_mulsc_mulb_yos113;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy113 = multm_reduce_mulsc_mulb_sq114 & multm_reduce_mulsc_mulb_yos114;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy114 = multm_reduce_mulsc_mulb_sq115 & multm_reduce_mulsc_mulb_yos115;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy115 = multm_reduce_mulsc_mulb_sq116 & multm_reduce_mulsc_mulb_yos116;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy116 = multm_reduce_mulsc_mulb_sq117 & multm_reduce_mulsc_mulb_yos117;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy117 = multm_reduce_mulsc_mulb_sq118 & multm_reduce_mulsc_mulb_yos118;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy118 = multm_reduce_mulsc_mulb_sq119 & multm_reduce_mulsc_mulb_yos119;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy119 = multm_reduce_mulsc_mulb_sq120 & multm_reduce_mulsc_mulb_yos120;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy120 = multm_reduce_mulsc_mulb_sq121 & multm_reduce_mulsc_mulb_yos121;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy121 = multm_reduce_mulsc_mulb_sq122 & multm_reduce_mulsc_mulb_yos122;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy122 = multm_reduce_mulsc_mulb_sq123 & multm_reduce_mulsc_mulb_yos123;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy123 = multm_reduce_mulsc_mulb_sq124 & multm_reduce_mulsc_mulb_yos124;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy124 = multm_reduce_mulsc_mulb_sq125 & multm_reduce_mulsc_mulb_yos125;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy125 = multm_reduce_mulsc_mulb_sq126 & multm_reduce_mulsc_mulb_yos126;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy126 = multm_reduce_mulsc_mulb_sq127 & multm_reduce_mulsc_mulb_yos127;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy127 = multm_reduce_mulsc_mulb_sq128 & multm_reduce_mulsc_mulb_yos128;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy128 = multm_reduce_mulsc_mulb_sq129 & multm_reduce_mulsc_mulb_yos129;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy129 = multm_reduce_mulsc_mulb_sq130 & multm_reduce_mulsc_mulb_yos130;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy130 = multm_reduce_mulsc_mulb_sq131 & multm_reduce_mulsc_mulb_yos131;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy131 = multm_reduce_mulsc_mulb_sq132 & multm_reduce_mulsc_mulb_yos132;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy132 = multm_reduce_mulsc_mulb_sq133 & multm_reduce_mulsc_mulb_yos133;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy133 = multm_reduce_mulsc_mulb_sq134 & multm_reduce_mulsc_mulb_yos134;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy134 = multm_reduce_mulsc_mulb_sq135 & multm_reduce_mulsc_mulb_yos135;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy135 = multm_reduce_mulsc_mulb_sq136 & multm_reduce_mulsc_mulb_yos136;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy136 = multm_reduce_mulsc_mulb_sq137 & multm_reduce_mulsc_mulb_yos137;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy137 = multm_reduce_mulsc_mulb_sq138 & multm_reduce_mulsc_mulb_yos138;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy138 = multm_reduce_mulsc_mulb_sq139 & multm_reduce_mulsc_mulb_yos139;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy139 = multm_reduce_mulsc_mulb_sq140 & multm_reduce_mulsc_mulb_yos140;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy140 = multm_reduce_mulsc_mulb_sq141 & multm_reduce_mulsc_mulb_yos141;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy141 = multm_reduce_mulsc_mulb_sq142 & multm_reduce_mulsc_mulb_yos142;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy142 = multm_reduce_mulsc_mulb_sq143 & multm_reduce_mulsc_mulb_yos143;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy143 = multm_reduce_mulsc_mulb_sq144 & multm_reduce_mulsc_mulb_yos144;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy144 = multm_reduce_mulsc_mulb_sq145 & multm_reduce_mulsc_mulb_yos145;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy145 = multm_reduce_mulsc_mulb_sq146 & multm_reduce_mulsc_mulb_yos146;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy146 = multm_reduce_mulsc_mulb_sq147 & multm_reduce_mulsc_mulb_yos147;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy147 = multm_reduce_mulsc_mulb_sq148 & multm_reduce_mulsc_mulb_yos148;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy148 = multm_reduce_mulsc_mulb_sq149 & multm_reduce_mulsc_mulb_yos149;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy149 = multm_reduce_mulsc_mulb_sq150 & multm_reduce_mulsc_mulb_yos150;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy150 = multm_reduce_mulsc_mulb_sq151 & multm_reduce_mulsc_mulb_yos151;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy151 = multm_reduce_mulsc_mulb_sq152 & multm_reduce_mulsc_mulb_yos152;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy152 = multm_reduce_mulsc_mulb_sq153 & multm_reduce_mulsc_mulb_yos153;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy153 = multm_reduce_mulsc_mulb_sq154 & multm_reduce_mulsc_mulb_yos154;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy154 = multm_reduce_mulsc_mulb_sq155 & multm_reduce_mulsc_mulb_yos155;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy155 = multm_reduce_mulsc_mulb_sq156 & multm_reduce_mulsc_mulb_yos156;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy156 = multm_reduce_mulsc_mulb_sq157 & multm_reduce_mulsc_mulb_yos157;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy157 = multm_reduce_mulsc_mulb_sq158 & multm_reduce_mulsc_mulb_yos158;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy158 = multm_reduce_mulsc_mulb_sq159 & multm_reduce_mulsc_mulb_yos159;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy159 = multm_reduce_mulsc_mulb_sq160 & multm_reduce_mulsc_mulb_yos160;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy160 = multm_reduce_mulsc_mulb_sq161 & multm_reduce_mulsc_mulb_yos161;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy161 = multm_reduce_mulsc_mulb_sq162 & multm_reduce_mulsc_mulb_yos162;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy162 = multm_reduce_mulsc_mulb_sq163 & multm_reduce_mulsc_mulb_yos163;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy163 = multm_reduce_mulsc_mulb_sq164 & multm_reduce_mulsc_mulb_yos164;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy164 = multm_reduce_mulsc_mulb_sq165 & multm_reduce_mulsc_mulb_yos165;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy165 = multm_reduce_mulsc_mulb_sq166 & multm_reduce_mulsc_mulb_yos166;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy166 = multm_reduce_mulsc_mulb_sq167 & multm_reduce_mulsc_mulb_yos167;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy167 = multm_reduce_mulsc_mulb_sq168 & multm_reduce_mulsc_mulb_yos168;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy168 = multm_reduce_mulsc_mulb_sq169 & multm_reduce_mulsc_mulb_yos169;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy169 = multm_reduce_mulsc_mulb_sq170 & multm_reduce_mulsc_mulb_yos170;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy170 = multm_reduce_mulsc_mulb_sq171 & multm_reduce_mulsc_mulb_yos171;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy171 = multm_reduce_mulsc_mulb_sq172 & multm_reduce_mulsc_mulb_yos172;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy172 = multm_reduce_mulsc_mulb_sq173 & multm_reduce_mulsc_mulb_yos173;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy173 = multm_reduce_mulsc_mulb_sq174 & multm_reduce_mulsc_mulb_yos174;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy174 = multm_reduce_mulsc_mulb_sq175 & multm_reduce_mulsc_mulb_yos175;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy175 = multm_reduce_mulsc_mulb_sq176 & multm_reduce_mulsc_mulb_yos176;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy176 = multm_reduce_mulsc_mulb_sq177 & multm_reduce_mulsc_mulb_yos177;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy177 = multm_reduce_mulsc_mulb_sq178 & multm_reduce_mulsc_mulb_yos178;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy178 = multm_reduce_mulsc_mulb_sq179 & multm_reduce_mulsc_mulb_yos179;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy179 = multm_reduce_mulsc_mulb_sq180 & multm_reduce_mulsc_mulb_yos180;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy180 = multm_reduce_mulsc_mulb_sq181 & multm_reduce_mulsc_mulb_yos181;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy181 = multm_reduce_mulsc_mulb_sq182 & multm_reduce_mulsc_mulb_yos182;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_wy182 = multm_reduce_mulsc_mulb_sq183 & multm_reduce_mulsc_mulb_yos183;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy0 = multm_reduce_mulsc_mulb_cq0 & multm_reduce_mulsc_mulb_yos1;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy1 = multm_reduce_mulsc_mulb_cq1 & multm_reduce_mulsc_mulb_yos2;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy2 = multm_reduce_mulsc_mulb_cq2 & multm_reduce_mulsc_mulb_yos3;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy3 = multm_reduce_mulsc_mulb_cq3 & multm_reduce_mulsc_mulb_yos4;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy4 = multm_reduce_mulsc_mulb_cq4 & multm_reduce_mulsc_mulb_yos5;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy5 = multm_reduce_mulsc_mulb_cq5 & multm_reduce_mulsc_mulb_yos6;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy6 = multm_reduce_mulsc_mulb_cq6 & multm_reduce_mulsc_mulb_yos7;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy7 = multm_reduce_mulsc_mulb_cq7 & multm_reduce_mulsc_mulb_yos8;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy8 = multm_reduce_mulsc_mulb_cq8 & multm_reduce_mulsc_mulb_yos9;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy9 = multm_reduce_mulsc_mulb_cq9 & multm_reduce_mulsc_mulb_yos10;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy10 = multm_reduce_mulsc_mulb_cq10 & multm_reduce_mulsc_mulb_yos11;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy11 = multm_reduce_mulsc_mulb_cq11 & multm_reduce_mulsc_mulb_yos12;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy12 = multm_reduce_mulsc_mulb_cq12 & multm_reduce_mulsc_mulb_yos13;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy13 = multm_reduce_mulsc_mulb_cq13 & multm_reduce_mulsc_mulb_yos14;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy14 = multm_reduce_mulsc_mulb_cq14 & multm_reduce_mulsc_mulb_yos15;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy15 = multm_reduce_mulsc_mulb_cq15 & multm_reduce_mulsc_mulb_yos16;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy16 = multm_reduce_mulsc_mulb_cq16 & multm_reduce_mulsc_mulb_yos17;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy17 = multm_reduce_mulsc_mulb_cq17 & multm_reduce_mulsc_mulb_yos18;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy18 = multm_reduce_mulsc_mulb_cq18 & multm_reduce_mulsc_mulb_yos19;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy19 = multm_reduce_mulsc_mulb_cq19 & multm_reduce_mulsc_mulb_yos20;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy20 = multm_reduce_mulsc_mulb_cq20 & multm_reduce_mulsc_mulb_yos21;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy21 = multm_reduce_mulsc_mulb_cq21 & multm_reduce_mulsc_mulb_yos22;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy22 = multm_reduce_mulsc_mulb_cq22 & multm_reduce_mulsc_mulb_yos23;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy23 = multm_reduce_mulsc_mulb_cq23 & multm_reduce_mulsc_mulb_yos24;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy24 = multm_reduce_mulsc_mulb_cq24 & multm_reduce_mulsc_mulb_yos25;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy25 = multm_reduce_mulsc_mulb_cq25 & multm_reduce_mulsc_mulb_yos26;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy26 = multm_reduce_mulsc_mulb_cq26 & multm_reduce_mulsc_mulb_yos27;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy27 = multm_reduce_mulsc_mulb_cq27 & multm_reduce_mulsc_mulb_yos28;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy28 = multm_reduce_mulsc_mulb_cq28 & multm_reduce_mulsc_mulb_yos29;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy29 = multm_reduce_mulsc_mulb_cq29 & multm_reduce_mulsc_mulb_yos30;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy30 = multm_reduce_mulsc_mulb_cq30 & multm_reduce_mulsc_mulb_yos31;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy31 = multm_reduce_mulsc_mulb_cq31 & multm_reduce_mulsc_mulb_yos32;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy32 = multm_reduce_mulsc_mulb_cq32 & multm_reduce_mulsc_mulb_yos33;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy33 = multm_reduce_mulsc_mulb_cq33 & multm_reduce_mulsc_mulb_yos34;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy34 = multm_reduce_mulsc_mulb_cq34 & multm_reduce_mulsc_mulb_yos35;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy35 = multm_reduce_mulsc_mulb_cq35 & multm_reduce_mulsc_mulb_yos36;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy36 = multm_reduce_mulsc_mulb_cq36 & multm_reduce_mulsc_mulb_yos37;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy37 = multm_reduce_mulsc_mulb_cq37 & multm_reduce_mulsc_mulb_yos38;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy38 = multm_reduce_mulsc_mulb_cq38 & multm_reduce_mulsc_mulb_yos39;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy39 = multm_reduce_mulsc_mulb_cq39 & multm_reduce_mulsc_mulb_yos40;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy40 = multm_reduce_mulsc_mulb_cq40 & multm_reduce_mulsc_mulb_yos41;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy41 = multm_reduce_mulsc_mulb_cq41 & multm_reduce_mulsc_mulb_yos42;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy42 = multm_reduce_mulsc_mulb_cq42 & multm_reduce_mulsc_mulb_yos43;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy43 = multm_reduce_mulsc_mulb_cq43 & multm_reduce_mulsc_mulb_yos44;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy44 = multm_reduce_mulsc_mulb_cq44 & multm_reduce_mulsc_mulb_yos45;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy45 = multm_reduce_mulsc_mulb_cq45 & multm_reduce_mulsc_mulb_yos46;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy46 = multm_reduce_mulsc_mulb_cq46 & multm_reduce_mulsc_mulb_yos47;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy47 = multm_reduce_mulsc_mulb_cq47 & multm_reduce_mulsc_mulb_yos48;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy48 = multm_reduce_mulsc_mulb_cq48 & multm_reduce_mulsc_mulb_yos49;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy49 = multm_reduce_mulsc_mulb_cq49 & multm_reduce_mulsc_mulb_yos50;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy50 = multm_reduce_mulsc_mulb_cq50 & multm_reduce_mulsc_mulb_yos51;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy51 = multm_reduce_mulsc_mulb_cq51 & multm_reduce_mulsc_mulb_yos52;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy52 = multm_reduce_mulsc_mulb_cq52 & multm_reduce_mulsc_mulb_yos53;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy53 = multm_reduce_mulsc_mulb_cq53 & multm_reduce_mulsc_mulb_yos54;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy54 = multm_reduce_mulsc_mulb_cq54 & multm_reduce_mulsc_mulb_yos55;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy55 = multm_reduce_mulsc_mulb_cq55 & multm_reduce_mulsc_mulb_yos56;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy56 = multm_reduce_mulsc_mulb_cq56 & multm_reduce_mulsc_mulb_yos57;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy57 = multm_reduce_mulsc_mulb_cq57 & multm_reduce_mulsc_mulb_yos58;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy58 = multm_reduce_mulsc_mulb_cq58 & multm_reduce_mulsc_mulb_yos59;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy59 = multm_reduce_mulsc_mulb_cq59 & multm_reduce_mulsc_mulb_yos60;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy60 = multm_reduce_mulsc_mulb_cq60 & multm_reduce_mulsc_mulb_yos61;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy61 = multm_reduce_mulsc_mulb_cq61 & multm_reduce_mulsc_mulb_yos62;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy62 = multm_reduce_mulsc_mulb_cq62 & multm_reduce_mulsc_mulb_yos63;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy63 = multm_reduce_mulsc_mulb_cq63 & multm_reduce_mulsc_mulb_yos64;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy64 = multm_reduce_mulsc_mulb_cq64 & multm_reduce_mulsc_mulb_yos65;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy65 = multm_reduce_mulsc_mulb_cq65 & multm_reduce_mulsc_mulb_yos66;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy66 = multm_reduce_mulsc_mulb_cq66 & multm_reduce_mulsc_mulb_yos67;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy67 = multm_reduce_mulsc_mulb_cq67 & multm_reduce_mulsc_mulb_yos68;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy68 = multm_reduce_mulsc_mulb_cq68 & multm_reduce_mulsc_mulb_yos69;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy69 = multm_reduce_mulsc_mulb_cq69 & multm_reduce_mulsc_mulb_yos70;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy70 = multm_reduce_mulsc_mulb_cq70 & multm_reduce_mulsc_mulb_yos71;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy71 = multm_reduce_mulsc_mulb_cq71 & multm_reduce_mulsc_mulb_yos72;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy72 = multm_reduce_mulsc_mulb_cq72 & multm_reduce_mulsc_mulb_yos73;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy73 = multm_reduce_mulsc_mulb_cq73 & multm_reduce_mulsc_mulb_yos74;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy74 = multm_reduce_mulsc_mulb_cq74 & multm_reduce_mulsc_mulb_yos75;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy75 = multm_reduce_mulsc_mulb_cq75 & multm_reduce_mulsc_mulb_yos76;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy76 = multm_reduce_mulsc_mulb_cq76 & multm_reduce_mulsc_mulb_yos77;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy77 = multm_reduce_mulsc_mulb_cq77 & multm_reduce_mulsc_mulb_yos78;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy78 = multm_reduce_mulsc_mulb_cq78 & multm_reduce_mulsc_mulb_yos79;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy79 = multm_reduce_mulsc_mulb_cq79 & multm_reduce_mulsc_mulb_yos80;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy80 = multm_reduce_mulsc_mulb_cq80 & multm_reduce_mulsc_mulb_yos81;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy81 = multm_reduce_mulsc_mulb_cq81 & multm_reduce_mulsc_mulb_yos82;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy82 = multm_reduce_mulsc_mulb_cq82 & multm_reduce_mulsc_mulb_yos83;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy83 = multm_reduce_mulsc_mulb_cq83 & multm_reduce_mulsc_mulb_yos84;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy84 = multm_reduce_mulsc_mulb_cq84 & multm_reduce_mulsc_mulb_yos85;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy85 = multm_reduce_mulsc_mulb_cq85 & multm_reduce_mulsc_mulb_yos86;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy86 = multm_reduce_mulsc_mulb_cq86 & multm_reduce_mulsc_mulb_yos87;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy87 = multm_reduce_mulsc_mulb_cq87 & multm_reduce_mulsc_mulb_yos88;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy88 = multm_reduce_mulsc_mulb_cq88 & multm_reduce_mulsc_mulb_yos89;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy89 = multm_reduce_mulsc_mulb_cq89 & multm_reduce_mulsc_mulb_yos90;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy90 = multm_reduce_mulsc_mulb_cq90 & multm_reduce_mulsc_mulb_yos91;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy91 = multm_reduce_mulsc_mulb_cq91 & multm_reduce_mulsc_mulb_yos92;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy92 = multm_reduce_mulsc_mulb_cq92 & multm_reduce_mulsc_mulb_yos93;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy93 = multm_reduce_mulsc_mulb_cq93 & multm_reduce_mulsc_mulb_yos94;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy94 = multm_reduce_mulsc_mulb_cq94 & multm_reduce_mulsc_mulb_yos95;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy95 = multm_reduce_mulsc_mulb_cq95 & multm_reduce_mulsc_mulb_yos96;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy96 = multm_reduce_mulsc_mulb_cq96 & multm_reduce_mulsc_mulb_yos97;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy97 = multm_reduce_mulsc_mulb_cq97 & multm_reduce_mulsc_mulb_yos98;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy98 = multm_reduce_mulsc_mulb_cq98 & multm_reduce_mulsc_mulb_yos99;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy99 = multm_reduce_mulsc_mulb_cq99 & multm_reduce_mulsc_mulb_yos100;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy100 = multm_reduce_mulsc_mulb_cq100 & multm_reduce_mulsc_mulb_yos101;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy101 = multm_reduce_mulsc_mulb_cq101 & multm_reduce_mulsc_mulb_yos102;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy102 = multm_reduce_mulsc_mulb_cq102 & multm_reduce_mulsc_mulb_yos103;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy103 = multm_reduce_mulsc_mulb_cq103 & multm_reduce_mulsc_mulb_yos104;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy104 = multm_reduce_mulsc_mulb_cq104 & multm_reduce_mulsc_mulb_yos105;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy105 = multm_reduce_mulsc_mulb_cq105 & multm_reduce_mulsc_mulb_yos106;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy106 = multm_reduce_mulsc_mulb_cq106 & multm_reduce_mulsc_mulb_yos107;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy107 = multm_reduce_mulsc_mulb_cq107 & multm_reduce_mulsc_mulb_yos108;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy108 = multm_reduce_mulsc_mulb_cq108 & multm_reduce_mulsc_mulb_yos109;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy109 = multm_reduce_mulsc_mulb_cq109 & multm_reduce_mulsc_mulb_yos110;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy110 = multm_reduce_mulsc_mulb_cq110 & multm_reduce_mulsc_mulb_yos111;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy111 = multm_reduce_mulsc_mulb_cq111 & multm_reduce_mulsc_mulb_yos112;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy112 = multm_reduce_mulsc_mulb_cq112 & multm_reduce_mulsc_mulb_yos113;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy113 = multm_reduce_mulsc_mulb_cq113 & multm_reduce_mulsc_mulb_yos114;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy114 = multm_reduce_mulsc_mulb_cq114 & multm_reduce_mulsc_mulb_yos115;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy115 = multm_reduce_mulsc_mulb_cq115 & multm_reduce_mulsc_mulb_yos116;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy116 = multm_reduce_mulsc_mulb_cq116 & multm_reduce_mulsc_mulb_yos117;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy117 = multm_reduce_mulsc_mulb_cq117 & multm_reduce_mulsc_mulb_yos118;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy118 = multm_reduce_mulsc_mulb_cq118 & multm_reduce_mulsc_mulb_yos119;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy119 = multm_reduce_mulsc_mulb_cq119 & multm_reduce_mulsc_mulb_yos120;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy120 = multm_reduce_mulsc_mulb_cq120 & multm_reduce_mulsc_mulb_yos121;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy121 = multm_reduce_mulsc_mulb_cq121 & multm_reduce_mulsc_mulb_yos122;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy122 = multm_reduce_mulsc_mulb_cq122 & multm_reduce_mulsc_mulb_yos123;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy123 = multm_reduce_mulsc_mulb_cq123 & multm_reduce_mulsc_mulb_yos124;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy124 = multm_reduce_mulsc_mulb_cq124 & multm_reduce_mulsc_mulb_yos125;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy125 = multm_reduce_mulsc_mulb_cq125 & multm_reduce_mulsc_mulb_yos126;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy126 = multm_reduce_mulsc_mulb_cq126 & multm_reduce_mulsc_mulb_yos127;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy127 = multm_reduce_mulsc_mulb_cq127 & multm_reduce_mulsc_mulb_yos128;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy128 = multm_reduce_mulsc_mulb_cq128 & multm_reduce_mulsc_mulb_yos129;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy129 = multm_reduce_mulsc_mulb_cq129 & multm_reduce_mulsc_mulb_yos130;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy130 = multm_reduce_mulsc_mulb_cq130 & multm_reduce_mulsc_mulb_yos131;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy131 = multm_reduce_mulsc_mulb_cq131 & multm_reduce_mulsc_mulb_yos132;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy132 = multm_reduce_mulsc_mulb_cq132 & multm_reduce_mulsc_mulb_yos133;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy133 = multm_reduce_mulsc_mulb_cq133 & multm_reduce_mulsc_mulb_yos134;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy134 = multm_reduce_mulsc_mulb_cq134 & multm_reduce_mulsc_mulb_yos135;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy135 = multm_reduce_mulsc_mulb_cq135 & multm_reduce_mulsc_mulb_yos136;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy136 = multm_reduce_mulsc_mulb_cq136 & multm_reduce_mulsc_mulb_yos137;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy137 = multm_reduce_mulsc_mulb_cq137 & multm_reduce_mulsc_mulb_yos138;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy138 = multm_reduce_mulsc_mulb_cq138 & multm_reduce_mulsc_mulb_yos139;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy139 = multm_reduce_mulsc_mulb_cq139 & multm_reduce_mulsc_mulb_yos140;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy140 = multm_reduce_mulsc_mulb_cq140 & multm_reduce_mulsc_mulb_yos141;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy141 = multm_reduce_mulsc_mulb_cq141 & multm_reduce_mulsc_mulb_yos142;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy142 = multm_reduce_mulsc_mulb_cq142 & multm_reduce_mulsc_mulb_yos143;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy143 = multm_reduce_mulsc_mulb_cq143 & multm_reduce_mulsc_mulb_yos144;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy144 = multm_reduce_mulsc_mulb_cq144 & multm_reduce_mulsc_mulb_yos145;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy145 = multm_reduce_mulsc_mulb_cq145 & multm_reduce_mulsc_mulb_yos146;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy146 = multm_reduce_mulsc_mulb_cq146 & multm_reduce_mulsc_mulb_yos147;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy147 = multm_reduce_mulsc_mulb_cq147 & multm_reduce_mulsc_mulb_yos148;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy148 = multm_reduce_mulsc_mulb_cq148 & multm_reduce_mulsc_mulb_yos149;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy149 = multm_reduce_mulsc_mulb_cq149 & multm_reduce_mulsc_mulb_yos150;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy150 = multm_reduce_mulsc_mulb_cq150 & multm_reduce_mulsc_mulb_yos151;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy151 = multm_reduce_mulsc_mulb_cq151 & multm_reduce_mulsc_mulb_yos152;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy152 = multm_reduce_mulsc_mulb_cq152 & multm_reduce_mulsc_mulb_yos153;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy153 = multm_reduce_mulsc_mulb_cq153 & multm_reduce_mulsc_mulb_yos154;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy154 = multm_reduce_mulsc_mulb_cq154 & multm_reduce_mulsc_mulb_yos155;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy155 = multm_reduce_mulsc_mulb_cq155 & multm_reduce_mulsc_mulb_yos156;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy156 = multm_reduce_mulsc_mulb_cq156 & multm_reduce_mulsc_mulb_yos157;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy157 = multm_reduce_mulsc_mulb_cq157 & multm_reduce_mulsc_mulb_yos158;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy158 = multm_reduce_mulsc_mulb_cq158 & multm_reduce_mulsc_mulb_yos159;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy159 = multm_reduce_mulsc_mulb_cq159 & multm_reduce_mulsc_mulb_yos160;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy160 = multm_reduce_mulsc_mulb_cq160 & multm_reduce_mulsc_mulb_yos161;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy161 = multm_reduce_mulsc_mulb_cq161 & multm_reduce_mulsc_mulb_yos162;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy162 = multm_reduce_mulsc_mulb_cq162 & multm_reduce_mulsc_mulb_yos163;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy163 = multm_reduce_mulsc_mulb_cq163 & multm_reduce_mulsc_mulb_yos164;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy164 = multm_reduce_mulsc_mulb_cq164 & multm_reduce_mulsc_mulb_yos165;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy165 = multm_reduce_mulsc_mulb_cq165 & multm_reduce_mulsc_mulb_yos166;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy166 = multm_reduce_mulsc_mulb_cq166 & multm_reduce_mulsc_mulb_yos167;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy167 = multm_reduce_mulsc_mulb_cq167 & multm_reduce_mulsc_mulb_yos168;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy168 = multm_reduce_mulsc_mulb_cq168 & multm_reduce_mulsc_mulb_yos169;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy169 = multm_reduce_mulsc_mulb_cq169 & multm_reduce_mulsc_mulb_yos170;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy170 = multm_reduce_mulsc_mulb_cq170 & multm_reduce_mulsc_mulb_yos171;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy171 = multm_reduce_mulsc_mulb_cq171 & multm_reduce_mulsc_mulb_yos172;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy172 = multm_reduce_mulsc_mulb_cq172 & multm_reduce_mulsc_mulb_yos173;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy173 = multm_reduce_mulsc_mulb_cq173 & multm_reduce_mulsc_mulb_yos174;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy174 = multm_reduce_mulsc_mulb_cq174 & multm_reduce_mulsc_mulb_yos175;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy175 = multm_reduce_mulsc_mulb_cq175 & multm_reduce_mulsc_mulb_yos176;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy176 = multm_reduce_mulsc_mulb_cq176 & multm_reduce_mulsc_mulb_yos177;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy177 = multm_reduce_mulsc_mulb_cq177 & multm_reduce_mulsc_mulb_yos178;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy178 = multm_reduce_mulsc_mulb_cq178 & multm_reduce_mulsc_mulb_yos179;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy179 = multm_reduce_mulsc_mulb_cq179 & multm_reduce_mulsc_mulb_yos180;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy180 = multm_reduce_mulsc_mulb_cq180 & multm_reduce_mulsc_mulb_yos181;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy181 = multm_reduce_mulsc_mulb_cq181 & multm_reduce_mulsc_mulb_yos182;
  assign multm_reduce_mulsc_mulb_add3b0_maj3b_xy182 = multm_reduce_mulsc_mulb_cq182 & multm_reduce_mulsc_mulb_yos183;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx0 = multm_reduce_mulsc_mulb_sq1 ^ multm_reduce_mulsc_mulb_cq0;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx1 = multm_reduce_mulsc_mulb_sq2 ^ multm_reduce_mulsc_mulb_cq1;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx2 = multm_reduce_mulsc_mulb_sq3 ^ multm_reduce_mulsc_mulb_cq2;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx3 = multm_reduce_mulsc_mulb_sq4 ^ multm_reduce_mulsc_mulb_cq3;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx4 = multm_reduce_mulsc_mulb_sq5 ^ multm_reduce_mulsc_mulb_cq4;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx5 = multm_reduce_mulsc_mulb_sq6 ^ multm_reduce_mulsc_mulb_cq5;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx6 = multm_reduce_mulsc_mulb_sq7 ^ multm_reduce_mulsc_mulb_cq6;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx7 = multm_reduce_mulsc_mulb_sq8 ^ multm_reduce_mulsc_mulb_cq7;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx8 = multm_reduce_mulsc_mulb_sq9 ^ multm_reduce_mulsc_mulb_cq8;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx9 = multm_reduce_mulsc_mulb_sq10 ^ multm_reduce_mulsc_mulb_cq9;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx10 = multm_reduce_mulsc_mulb_sq11 ^ multm_reduce_mulsc_mulb_cq10;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx11 = multm_reduce_mulsc_mulb_sq12 ^ multm_reduce_mulsc_mulb_cq11;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx12 = multm_reduce_mulsc_mulb_sq13 ^ multm_reduce_mulsc_mulb_cq12;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx13 = multm_reduce_mulsc_mulb_sq14 ^ multm_reduce_mulsc_mulb_cq13;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx14 = multm_reduce_mulsc_mulb_sq15 ^ multm_reduce_mulsc_mulb_cq14;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx15 = multm_reduce_mulsc_mulb_sq16 ^ multm_reduce_mulsc_mulb_cq15;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx16 = multm_reduce_mulsc_mulb_sq17 ^ multm_reduce_mulsc_mulb_cq16;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx17 = multm_reduce_mulsc_mulb_sq18 ^ multm_reduce_mulsc_mulb_cq17;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx18 = multm_reduce_mulsc_mulb_sq19 ^ multm_reduce_mulsc_mulb_cq18;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx19 = multm_reduce_mulsc_mulb_sq20 ^ multm_reduce_mulsc_mulb_cq19;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx20 = multm_reduce_mulsc_mulb_sq21 ^ multm_reduce_mulsc_mulb_cq20;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx21 = multm_reduce_mulsc_mulb_sq22 ^ multm_reduce_mulsc_mulb_cq21;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx22 = multm_reduce_mulsc_mulb_sq23 ^ multm_reduce_mulsc_mulb_cq22;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx23 = multm_reduce_mulsc_mulb_sq24 ^ multm_reduce_mulsc_mulb_cq23;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx24 = multm_reduce_mulsc_mulb_sq25 ^ multm_reduce_mulsc_mulb_cq24;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx25 = multm_reduce_mulsc_mulb_sq26 ^ multm_reduce_mulsc_mulb_cq25;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx26 = multm_reduce_mulsc_mulb_sq27 ^ multm_reduce_mulsc_mulb_cq26;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx27 = multm_reduce_mulsc_mulb_sq28 ^ multm_reduce_mulsc_mulb_cq27;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx28 = multm_reduce_mulsc_mulb_sq29 ^ multm_reduce_mulsc_mulb_cq28;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx29 = multm_reduce_mulsc_mulb_sq30 ^ multm_reduce_mulsc_mulb_cq29;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx30 = multm_reduce_mulsc_mulb_sq31 ^ multm_reduce_mulsc_mulb_cq30;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx31 = multm_reduce_mulsc_mulb_sq32 ^ multm_reduce_mulsc_mulb_cq31;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx32 = multm_reduce_mulsc_mulb_sq33 ^ multm_reduce_mulsc_mulb_cq32;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx33 = multm_reduce_mulsc_mulb_sq34 ^ multm_reduce_mulsc_mulb_cq33;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx34 = multm_reduce_mulsc_mulb_sq35 ^ multm_reduce_mulsc_mulb_cq34;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx35 = multm_reduce_mulsc_mulb_sq36 ^ multm_reduce_mulsc_mulb_cq35;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx36 = multm_reduce_mulsc_mulb_sq37 ^ multm_reduce_mulsc_mulb_cq36;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx37 = multm_reduce_mulsc_mulb_sq38 ^ multm_reduce_mulsc_mulb_cq37;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx38 = multm_reduce_mulsc_mulb_sq39 ^ multm_reduce_mulsc_mulb_cq38;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx39 = multm_reduce_mulsc_mulb_sq40 ^ multm_reduce_mulsc_mulb_cq39;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx40 = multm_reduce_mulsc_mulb_sq41 ^ multm_reduce_mulsc_mulb_cq40;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx41 = multm_reduce_mulsc_mulb_sq42 ^ multm_reduce_mulsc_mulb_cq41;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx42 = multm_reduce_mulsc_mulb_sq43 ^ multm_reduce_mulsc_mulb_cq42;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx43 = multm_reduce_mulsc_mulb_sq44 ^ multm_reduce_mulsc_mulb_cq43;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx44 = multm_reduce_mulsc_mulb_sq45 ^ multm_reduce_mulsc_mulb_cq44;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx45 = multm_reduce_mulsc_mulb_sq46 ^ multm_reduce_mulsc_mulb_cq45;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx46 = multm_reduce_mulsc_mulb_sq47 ^ multm_reduce_mulsc_mulb_cq46;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx47 = multm_reduce_mulsc_mulb_sq48 ^ multm_reduce_mulsc_mulb_cq47;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx48 = multm_reduce_mulsc_mulb_sq49 ^ multm_reduce_mulsc_mulb_cq48;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx49 = multm_reduce_mulsc_mulb_sq50 ^ multm_reduce_mulsc_mulb_cq49;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx50 = multm_reduce_mulsc_mulb_sq51 ^ multm_reduce_mulsc_mulb_cq50;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx51 = multm_reduce_mulsc_mulb_sq52 ^ multm_reduce_mulsc_mulb_cq51;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx52 = multm_reduce_mulsc_mulb_sq53 ^ multm_reduce_mulsc_mulb_cq52;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx53 = multm_reduce_mulsc_mulb_sq54 ^ multm_reduce_mulsc_mulb_cq53;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx54 = multm_reduce_mulsc_mulb_sq55 ^ multm_reduce_mulsc_mulb_cq54;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx55 = multm_reduce_mulsc_mulb_sq56 ^ multm_reduce_mulsc_mulb_cq55;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx56 = multm_reduce_mulsc_mulb_sq57 ^ multm_reduce_mulsc_mulb_cq56;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx57 = multm_reduce_mulsc_mulb_sq58 ^ multm_reduce_mulsc_mulb_cq57;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx58 = multm_reduce_mulsc_mulb_sq59 ^ multm_reduce_mulsc_mulb_cq58;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx59 = multm_reduce_mulsc_mulb_sq60 ^ multm_reduce_mulsc_mulb_cq59;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx60 = multm_reduce_mulsc_mulb_sq61 ^ multm_reduce_mulsc_mulb_cq60;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx61 = multm_reduce_mulsc_mulb_sq62 ^ multm_reduce_mulsc_mulb_cq61;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx62 = multm_reduce_mulsc_mulb_sq63 ^ multm_reduce_mulsc_mulb_cq62;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx63 = multm_reduce_mulsc_mulb_sq64 ^ multm_reduce_mulsc_mulb_cq63;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx64 = multm_reduce_mulsc_mulb_sq65 ^ multm_reduce_mulsc_mulb_cq64;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx65 = multm_reduce_mulsc_mulb_sq66 ^ multm_reduce_mulsc_mulb_cq65;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx66 = multm_reduce_mulsc_mulb_sq67 ^ multm_reduce_mulsc_mulb_cq66;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx67 = multm_reduce_mulsc_mulb_sq68 ^ multm_reduce_mulsc_mulb_cq67;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx68 = multm_reduce_mulsc_mulb_sq69 ^ multm_reduce_mulsc_mulb_cq68;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx69 = multm_reduce_mulsc_mulb_sq70 ^ multm_reduce_mulsc_mulb_cq69;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx70 = multm_reduce_mulsc_mulb_sq71 ^ multm_reduce_mulsc_mulb_cq70;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx71 = multm_reduce_mulsc_mulb_sq72 ^ multm_reduce_mulsc_mulb_cq71;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx72 = multm_reduce_mulsc_mulb_sq73 ^ multm_reduce_mulsc_mulb_cq72;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx73 = multm_reduce_mulsc_mulb_sq74 ^ multm_reduce_mulsc_mulb_cq73;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx74 = multm_reduce_mulsc_mulb_sq75 ^ multm_reduce_mulsc_mulb_cq74;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx75 = multm_reduce_mulsc_mulb_sq76 ^ multm_reduce_mulsc_mulb_cq75;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx76 = multm_reduce_mulsc_mulb_sq77 ^ multm_reduce_mulsc_mulb_cq76;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx77 = multm_reduce_mulsc_mulb_sq78 ^ multm_reduce_mulsc_mulb_cq77;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx78 = multm_reduce_mulsc_mulb_sq79 ^ multm_reduce_mulsc_mulb_cq78;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx79 = multm_reduce_mulsc_mulb_sq80 ^ multm_reduce_mulsc_mulb_cq79;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx80 = multm_reduce_mulsc_mulb_sq81 ^ multm_reduce_mulsc_mulb_cq80;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx81 = multm_reduce_mulsc_mulb_sq82 ^ multm_reduce_mulsc_mulb_cq81;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx82 = multm_reduce_mulsc_mulb_sq83 ^ multm_reduce_mulsc_mulb_cq82;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx83 = multm_reduce_mulsc_mulb_sq84 ^ multm_reduce_mulsc_mulb_cq83;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx84 = multm_reduce_mulsc_mulb_sq85 ^ multm_reduce_mulsc_mulb_cq84;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx85 = multm_reduce_mulsc_mulb_sq86 ^ multm_reduce_mulsc_mulb_cq85;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx86 = multm_reduce_mulsc_mulb_sq87 ^ multm_reduce_mulsc_mulb_cq86;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx87 = multm_reduce_mulsc_mulb_sq88 ^ multm_reduce_mulsc_mulb_cq87;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx88 = multm_reduce_mulsc_mulb_sq89 ^ multm_reduce_mulsc_mulb_cq88;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx89 = multm_reduce_mulsc_mulb_sq90 ^ multm_reduce_mulsc_mulb_cq89;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx90 = multm_reduce_mulsc_mulb_sq91 ^ multm_reduce_mulsc_mulb_cq90;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx91 = multm_reduce_mulsc_mulb_sq92 ^ multm_reduce_mulsc_mulb_cq91;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx92 = multm_reduce_mulsc_mulb_sq93 ^ multm_reduce_mulsc_mulb_cq92;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx93 = multm_reduce_mulsc_mulb_sq94 ^ multm_reduce_mulsc_mulb_cq93;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx94 = multm_reduce_mulsc_mulb_sq95 ^ multm_reduce_mulsc_mulb_cq94;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx95 = multm_reduce_mulsc_mulb_sq96 ^ multm_reduce_mulsc_mulb_cq95;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx96 = multm_reduce_mulsc_mulb_sq97 ^ multm_reduce_mulsc_mulb_cq96;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx97 = multm_reduce_mulsc_mulb_sq98 ^ multm_reduce_mulsc_mulb_cq97;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx98 = multm_reduce_mulsc_mulb_sq99 ^ multm_reduce_mulsc_mulb_cq98;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx99 = multm_reduce_mulsc_mulb_sq100 ^ multm_reduce_mulsc_mulb_cq99;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx100 = multm_reduce_mulsc_mulb_sq101 ^ multm_reduce_mulsc_mulb_cq100;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx101 = multm_reduce_mulsc_mulb_sq102 ^ multm_reduce_mulsc_mulb_cq101;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx102 = multm_reduce_mulsc_mulb_sq103 ^ multm_reduce_mulsc_mulb_cq102;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx103 = multm_reduce_mulsc_mulb_sq104 ^ multm_reduce_mulsc_mulb_cq103;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx104 = multm_reduce_mulsc_mulb_sq105 ^ multm_reduce_mulsc_mulb_cq104;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx105 = multm_reduce_mulsc_mulb_sq106 ^ multm_reduce_mulsc_mulb_cq105;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx106 = multm_reduce_mulsc_mulb_sq107 ^ multm_reduce_mulsc_mulb_cq106;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx107 = multm_reduce_mulsc_mulb_sq108 ^ multm_reduce_mulsc_mulb_cq107;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx108 = multm_reduce_mulsc_mulb_sq109 ^ multm_reduce_mulsc_mulb_cq108;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx109 = multm_reduce_mulsc_mulb_sq110 ^ multm_reduce_mulsc_mulb_cq109;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx110 = multm_reduce_mulsc_mulb_sq111 ^ multm_reduce_mulsc_mulb_cq110;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx111 = multm_reduce_mulsc_mulb_sq112 ^ multm_reduce_mulsc_mulb_cq111;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx112 = multm_reduce_mulsc_mulb_sq113 ^ multm_reduce_mulsc_mulb_cq112;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx113 = multm_reduce_mulsc_mulb_sq114 ^ multm_reduce_mulsc_mulb_cq113;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx114 = multm_reduce_mulsc_mulb_sq115 ^ multm_reduce_mulsc_mulb_cq114;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx115 = multm_reduce_mulsc_mulb_sq116 ^ multm_reduce_mulsc_mulb_cq115;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx116 = multm_reduce_mulsc_mulb_sq117 ^ multm_reduce_mulsc_mulb_cq116;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx117 = multm_reduce_mulsc_mulb_sq118 ^ multm_reduce_mulsc_mulb_cq117;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx118 = multm_reduce_mulsc_mulb_sq119 ^ multm_reduce_mulsc_mulb_cq118;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx119 = multm_reduce_mulsc_mulb_sq120 ^ multm_reduce_mulsc_mulb_cq119;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx120 = multm_reduce_mulsc_mulb_sq121 ^ multm_reduce_mulsc_mulb_cq120;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx121 = multm_reduce_mulsc_mulb_sq122 ^ multm_reduce_mulsc_mulb_cq121;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx122 = multm_reduce_mulsc_mulb_sq123 ^ multm_reduce_mulsc_mulb_cq122;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx123 = multm_reduce_mulsc_mulb_sq124 ^ multm_reduce_mulsc_mulb_cq123;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx124 = multm_reduce_mulsc_mulb_sq125 ^ multm_reduce_mulsc_mulb_cq124;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx125 = multm_reduce_mulsc_mulb_sq126 ^ multm_reduce_mulsc_mulb_cq125;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx126 = multm_reduce_mulsc_mulb_sq127 ^ multm_reduce_mulsc_mulb_cq126;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx127 = multm_reduce_mulsc_mulb_sq128 ^ multm_reduce_mulsc_mulb_cq127;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx128 = multm_reduce_mulsc_mulb_sq129 ^ multm_reduce_mulsc_mulb_cq128;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx129 = multm_reduce_mulsc_mulb_sq130 ^ multm_reduce_mulsc_mulb_cq129;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx130 = multm_reduce_mulsc_mulb_sq131 ^ multm_reduce_mulsc_mulb_cq130;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx131 = multm_reduce_mulsc_mulb_sq132 ^ multm_reduce_mulsc_mulb_cq131;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx132 = multm_reduce_mulsc_mulb_sq133 ^ multm_reduce_mulsc_mulb_cq132;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx133 = multm_reduce_mulsc_mulb_sq134 ^ multm_reduce_mulsc_mulb_cq133;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx134 = multm_reduce_mulsc_mulb_sq135 ^ multm_reduce_mulsc_mulb_cq134;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx135 = multm_reduce_mulsc_mulb_sq136 ^ multm_reduce_mulsc_mulb_cq135;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx136 = multm_reduce_mulsc_mulb_sq137 ^ multm_reduce_mulsc_mulb_cq136;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx137 = multm_reduce_mulsc_mulb_sq138 ^ multm_reduce_mulsc_mulb_cq137;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx138 = multm_reduce_mulsc_mulb_sq139 ^ multm_reduce_mulsc_mulb_cq138;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx139 = multm_reduce_mulsc_mulb_sq140 ^ multm_reduce_mulsc_mulb_cq139;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx140 = multm_reduce_mulsc_mulb_sq141 ^ multm_reduce_mulsc_mulb_cq140;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx141 = multm_reduce_mulsc_mulb_sq142 ^ multm_reduce_mulsc_mulb_cq141;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx142 = multm_reduce_mulsc_mulb_sq143 ^ multm_reduce_mulsc_mulb_cq142;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx143 = multm_reduce_mulsc_mulb_sq144 ^ multm_reduce_mulsc_mulb_cq143;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx144 = multm_reduce_mulsc_mulb_sq145 ^ multm_reduce_mulsc_mulb_cq144;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx145 = multm_reduce_mulsc_mulb_sq146 ^ multm_reduce_mulsc_mulb_cq145;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx146 = multm_reduce_mulsc_mulb_sq147 ^ multm_reduce_mulsc_mulb_cq146;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx147 = multm_reduce_mulsc_mulb_sq148 ^ multm_reduce_mulsc_mulb_cq147;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx148 = multm_reduce_mulsc_mulb_sq149 ^ multm_reduce_mulsc_mulb_cq148;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx149 = multm_reduce_mulsc_mulb_sq150 ^ multm_reduce_mulsc_mulb_cq149;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx150 = multm_reduce_mulsc_mulb_sq151 ^ multm_reduce_mulsc_mulb_cq150;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx151 = multm_reduce_mulsc_mulb_sq152 ^ multm_reduce_mulsc_mulb_cq151;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx152 = multm_reduce_mulsc_mulb_sq153 ^ multm_reduce_mulsc_mulb_cq152;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx153 = multm_reduce_mulsc_mulb_sq154 ^ multm_reduce_mulsc_mulb_cq153;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx154 = multm_reduce_mulsc_mulb_sq155 ^ multm_reduce_mulsc_mulb_cq154;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx155 = multm_reduce_mulsc_mulb_sq156 ^ multm_reduce_mulsc_mulb_cq155;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx156 = multm_reduce_mulsc_mulb_sq157 ^ multm_reduce_mulsc_mulb_cq156;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx157 = multm_reduce_mulsc_mulb_sq158 ^ multm_reduce_mulsc_mulb_cq157;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx158 = multm_reduce_mulsc_mulb_sq159 ^ multm_reduce_mulsc_mulb_cq158;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx159 = multm_reduce_mulsc_mulb_sq160 ^ multm_reduce_mulsc_mulb_cq159;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx160 = multm_reduce_mulsc_mulb_sq161 ^ multm_reduce_mulsc_mulb_cq160;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx161 = multm_reduce_mulsc_mulb_sq162 ^ multm_reduce_mulsc_mulb_cq161;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx162 = multm_reduce_mulsc_mulb_sq163 ^ multm_reduce_mulsc_mulb_cq162;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx163 = multm_reduce_mulsc_mulb_sq164 ^ multm_reduce_mulsc_mulb_cq163;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx164 = multm_reduce_mulsc_mulb_sq165 ^ multm_reduce_mulsc_mulb_cq164;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx165 = multm_reduce_mulsc_mulb_sq166 ^ multm_reduce_mulsc_mulb_cq165;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx166 = multm_reduce_mulsc_mulb_sq167 ^ multm_reduce_mulsc_mulb_cq166;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx167 = multm_reduce_mulsc_mulb_sq168 ^ multm_reduce_mulsc_mulb_cq167;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx168 = multm_reduce_mulsc_mulb_sq169 ^ multm_reduce_mulsc_mulb_cq168;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx169 = multm_reduce_mulsc_mulb_sq170 ^ multm_reduce_mulsc_mulb_cq169;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx170 = multm_reduce_mulsc_mulb_sq171 ^ multm_reduce_mulsc_mulb_cq170;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx171 = multm_reduce_mulsc_mulb_sq172 ^ multm_reduce_mulsc_mulb_cq171;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx172 = multm_reduce_mulsc_mulb_sq173 ^ multm_reduce_mulsc_mulb_cq172;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx173 = multm_reduce_mulsc_mulb_sq174 ^ multm_reduce_mulsc_mulb_cq173;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx174 = multm_reduce_mulsc_mulb_sq175 ^ multm_reduce_mulsc_mulb_cq174;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx175 = multm_reduce_mulsc_mulb_sq176 ^ multm_reduce_mulsc_mulb_cq175;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx176 = multm_reduce_mulsc_mulb_sq177 ^ multm_reduce_mulsc_mulb_cq176;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx177 = multm_reduce_mulsc_mulb_sq178 ^ multm_reduce_mulsc_mulb_cq177;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx178 = multm_reduce_mulsc_mulb_sq179 ^ multm_reduce_mulsc_mulb_cq178;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx179 = multm_reduce_mulsc_mulb_sq180 ^ multm_reduce_mulsc_mulb_cq179;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx180 = multm_reduce_mulsc_mulb_sq181 ^ multm_reduce_mulsc_mulb_cq180;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx181 = multm_reduce_mulsc_mulb_sq182 ^ multm_reduce_mulsc_mulb_cq181;
  assign multm_reduce_mulsc_mulb_add3b0_xor3b_wx182 = multm_reduce_mulsc_mulb_sq183 ^ multm_reduce_mulsc_mulb_cq182;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx0 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx0 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy0;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx1 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx1 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy1;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx2 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx2 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy2;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx3 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx3 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy3;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx4 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx4 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy4;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx5 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx5 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy5;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx6 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx6 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy6;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx7 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx7 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy7;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx8 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx8 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy8;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx9 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx9 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy9;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx10 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx10 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy10;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx11 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx11 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy11;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx12 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx12 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy12;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx13 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx13 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy13;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx14 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx14 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy14;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx15 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx15 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy15;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx16 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx16 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy16;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx17 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx17 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy17;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx18 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx18 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy18;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx19 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx19 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy19;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx20 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx20 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy20;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx21 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx21 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy21;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx22 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx22 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy22;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx23 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx23 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy23;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx24 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx24 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy24;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx25 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx25 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy25;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx26 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx26 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy26;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx27 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx27 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy27;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx28 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx28 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy28;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx29 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx29 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy29;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx30 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx30 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy30;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx31 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx31 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy31;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx32 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx32 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy32;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx33 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx33 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy33;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx34 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx34 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy34;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx35 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx35 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy35;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx36 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx36 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy36;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx37 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx37 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy37;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx38 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx38 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy38;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx39 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx39 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy39;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx40 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx40 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy40;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx41 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx41 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy41;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx42 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx42 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy42;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx43 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx43 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy43;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx44 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx44 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy44;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx45 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx45 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy45;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx46 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx46 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy46;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx47 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx47 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy47;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx48 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx48 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy48;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx49 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx49 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy49;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx50 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx50 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy50;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx51 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx51 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy51;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx52 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx52 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy52;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx53 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx53 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy53;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx54 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx54 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy54;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx55 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx55 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy55;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx56 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx56 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy56;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx57 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx57 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy57;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx58 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx58 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy58;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx59 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx59 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy59;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx60 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx60 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy60;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx61 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx61 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy61;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx62 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx62 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy62;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx63 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx63 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy63;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx64 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx64 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy64;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx65 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx65 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy65;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx66 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx66 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy66;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx67 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx67 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy67;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx68 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx68 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy68;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx69 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx69 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy69;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx70 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx70 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy70;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx71 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx71 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy71;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx72 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx72 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy72;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx73 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx73 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy73;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx74 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx74 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy74;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx75 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx75 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy75;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx76 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx76 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy76;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx77 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx77 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy77;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx78 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx78 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy78;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx79 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx79 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy79;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx80 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx80 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy80;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx81 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx81 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy81;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx82 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx82 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy82;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx83 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx83 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy83;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx84 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx84 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy84;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx85 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx85 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy85;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx86 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx86 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy86;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx87 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx87 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy87;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx88 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx88 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy88;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx89 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx89 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy89;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx90 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx90 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy90;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx91 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx91 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy91;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx92 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx92 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy92;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx93 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx93 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy93;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx94 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx94 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy94;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx95 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx95 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy95;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx96 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx96 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy96;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx97 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx97 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy97;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx98 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx98 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy98;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx99 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx99 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy99;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx100 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx100 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy100;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx101 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx101 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy101;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx102 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx102 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy102;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx103 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx103 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy103;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx104 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx104 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy104;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx105 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx105 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy105;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx106 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx106 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy106;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx107 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx107 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy107;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx108 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx108 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy108;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx109 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx109 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy109;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx110 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx110 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy110;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx111 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx111 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy111;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx112 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx112 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy112;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx113 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx113 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy113;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx114 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx114 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy114;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx115 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx115 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy115;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx116 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx116 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy116;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx117 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx117 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy117;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx118 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx118 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy118;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx119 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx119 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy119;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx120 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx120 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy120;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx121 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx121 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy121;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx122 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx122 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy122;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx123 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx123 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy123;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx124 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx124 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy124;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx125 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx125 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy125;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx126 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx126 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy126;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx127 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx127 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy127;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx128 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx128 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy128;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx129 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx129 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy129;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx130 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx130 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy130;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx131 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx131 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy131;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx132 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx132 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy132;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx133 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx133 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy133;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx134 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx134 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy134;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx135 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx135 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy135;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx136 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx136 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy136;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx137 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx137 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy137;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx138 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx138 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy138;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx139 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx139 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy139;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx140 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx140 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy140;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx141 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx141 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy141;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx142 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx142 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy142;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx143 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx143 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy143;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx144 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx144 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy144;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx145 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx145 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy145;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx146 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx146 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy146;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx147 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx147 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy147;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx148 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx148 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy148;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx149 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx149 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy149;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx150 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx150 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy150;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx151 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx151 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy151;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx152 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx152 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy152;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx153 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx153 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy153;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx154 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx154 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy154;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx155 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx155 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy155;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx156 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx156 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy156;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx157 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx157 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy157;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx158 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx158 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy158;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx159 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx159 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy159;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx160 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx160 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy160;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx161 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx161 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy161;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx162 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx162 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy162;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx163 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx163 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy163;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx164 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx164 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy164;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx165 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx165 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy165;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx166 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx166 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy166;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx167 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx167 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy167;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx168 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx168 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy168;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx169 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx169 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy169;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx170 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx170 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy170;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx171 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx171 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy171;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx172 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx172 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy172;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx173 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx173 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy173;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx174 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx174 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy174;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx175 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx175 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy175;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx176 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx176 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy176;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx177 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx177 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy177;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx178 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx178 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy178;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx179 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx179 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy179;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx180 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx180 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy180;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx181 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx181 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy181;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx182 = multm_reduce_mulsc_mulb_add3b1_maj3b_wx182 | multm_reduce_mulsc_mulb_add3b1_maj3b_wy182;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx0 = multm_reduce_mulsc_mulb_yoc0 & multm_reduce_mulsc_mulb_ps0;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx1 = multm_reduce_mulsc_mulb_yoc1 & multm_reduce_mulsc_mulb_ps1;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx2 = multm_reduce_mulsc_mulb_yoc2 & multm_reduce_mulsc_mulb_ps2;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx3 = multm_reduce_mulsc_mulb_yoc3 & multm_reduce_mulsc_mulb_ps3;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx4 = multm_reduce_mulsc_mulb_yoc4 & multm_reduce_mulsc_mulb_ps4;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx5 = multm_reduce_mulsc_mulb_yoc5 & multm_reduce_mulsc_mulb_ps5;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx6 = multm_reduce_mulsc_mulb_yoc6 & multm_reduce_mulsc_mulb_ps6;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx7 = multm_reduce_mulsc_mulb_yoc7 & multm_reduce_mulsc_mulb_ps7;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx8 = multm_reduce_mulsc_mulb_yoc8 & multm_reduce_mulsc_mulb_ps8;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx9 = multm_reduce_mulsc_mulb_yoc9 & multm_reduce_mulsc_mulb_ps9;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx10 = multm_reduce_mulsc_mulb_yoc10 & multm_reduce_mulsc_mulb_ps10;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx11 = multm_reduce_mulsc_mulb_yoc11 & multm_reduce_mulsc_mulb_ps11;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx12 = multm_reduce_mulsc_mulb_yoc12 & multm_reduce_mulsc_mulb_ps12;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx13 = multm_reduce_mulsc_mulb_yoc13 & multm_reduce_mulsc_mulb_ps13;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx14 = multm_reduce_mulsc_mulb_yoc14 & multm_reduce_mulsc_mulb_ps14;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx15 = multm_reduce_mulsc_mulb_yoc15 & multm_reduce_mulsc_mulb_ps15;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx16 = multm_reduce_mulsc_mulb_yoc16 & multm_reduce_mulsc_mulb_ps16;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx17 = multm_reduce_mulsc_mulb_yoc17 & multm_reduce_mulsc_mulb_ps17;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx18 = multm_reduce_mulsc_mulb_yoc18 & multm_reduce_mulsc_mulb_ps18;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx19 = multm_reduce_mulsc_mulb_yoc19 & multm_reduce_mulsc_mulb_ps19;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx20 = multm_reduce_mulsc_mulb_yoc20 & multm_reduce_mulsc_mulb_ps20;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx21 = multm_reduce_mulsc_mulb_yoc21 & multm_reduce_mulsc_mulb_ps21;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx22 = multm_reduce_mulsc_mulb_yoc22 & multm_reduce_mulsc_mulb_ps22;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx23 = multm_reduce_mulsc_mulb_yoc23 & multm_reduce_mulsc_mulb_ps23;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx24 = multm_reduce_mulsc_mulb_yoc24 & multm_reduce_mulsc_mulb_ps24;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx25 = multm_reduce_mulsc_mulb_yoc25 & multm_reduce_mulsc_mulb_ps25;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx26 = multm_reduce_mulsc_mulb_yoc26 & multm_reduce_mulsc_mulb_ps26;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx27 = multm_reduce_mulsc_mulb_yoc27 & multm_reduce_mulsc_mulb_ps27;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx28 = multm_reduce_mulsc_mulb_yoc28 & multm_reduce_mulsc_mulb_ps28;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx29 = multm_reduce_mulsc_mulb_yoc29 & multm_reduce_mulsc_mulb_ps29;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx30 = multm_reduce_mulsc_mulb_yoc30 & multm_reduce_mulsc_mulb_ps30;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx31 = multm_reduce_mulsc_mulb_yoc31 & multm_reduce_mulsc_mulb_ps31;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx32 = multm_reduce_mulsc_mulb_yoc32 & multm_reduce_mulsc_mulb_ps32;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx33 = multm_reduce_mulsc_mulb_yoc33 & multm_reduce_mulsc_mulb_ps33;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx34 = multm_reduce_mulsc_mulb_yoc34 & multm_reduce_mulsc_mulb_ps34;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx35 = multm_reduce_mulsc_mulb_yoc35 & multm_reduce_mulsc_mulb_ps35;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx36 = multm_reduce_mulsc_mulb_yoc36 & multm_reduce_mulsc_mulb_ps36;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx37 = multm_reduce_mulsc_mulb_yoc37 & multm_reduce_mulsc_mulb_ps37;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx38 = multm_reduce_mulsc_mulb_yoc38 & multm_reduce_mulsc_mulb_ps38;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx39 = multm_reduce_mulsc_mulb_yoc39 & multm_reduce_mulsc_mulb_ps39;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx40 = multm_reduce_mulsc_mulb_yoc40 & multm_reduce_mulsc_mulb_ps40;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx41 = multm_reduce_mulsc_mulb_yoc41 & multm_reduce_mulsc_mulb_ps41;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx42 = multm_reduce_mulsc_mulb_yoc42 & multm_reduce_mulsc_mulb_ps42;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx43 = multm_reduce_mulsc_mulb_yoc43 & multm_reduce_mulsc_mulb_ps43;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx44 = multm_reduce_mulsc_mulb_yoc44 & multm_reduce_mulsc_mulb_ps44;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx45 = multm_reduce_mulsc_mulb_yoc45 & multm_reduce_mulsc_mulb_ps45;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx46 = multm_reduce_mulsc_mulb_yoc46 & multm_reduce_mulsc_mulb_ps46;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx47 = multm_reduce_mulsc_mulb_yoc47 & multm_reduce_mulsc_mulb_ps47;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx48 = multm_reduce_mulsc_mulb_yoc48 & multm_reduce_mulsc_mulb_ps48;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx49 = multm_reduce_mulsc_mulb_yoc49 & multm_reduce_mulsc_mulb_ps49;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx50 = multm_reduce_mulsc_mulb_yoc50 & multm_reduce_mulsc_mulb_ps50;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx51 = multm_reduce_mulsc_mulb_yoc51 & multm_reduce_mulsc_mulb_ps51;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx52 = multm_reduce_mulsc_mulb_yoc52 & multm_reduce_mulsc_mulb_ps52;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx53 = multm_reduce_mulsc_mulb_yoc53 & multm_reduce_mulsc_mulb_ps53;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx54 = multm_reduce_mulsc_mulb_yoc54 & multm_reduce_mulsc_mulb_ps54;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx55 = multm_reduce_mulsc_mulb_yoc55 & multm_reduce_mulsc_mulb_ps55;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx56 = multm_reduce_mulsc_mulb_yoc56 & multm_reduce_mulsc_mulb_ps56;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx57 = multm_reduce_mulsc_mulb_yoc57 & multm_reduce_mulsc_mulb_ps57;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx58 = multm_reduce_mulsc_mulb_yoc58 & multm_reduce_mulsc_mulb_ps58;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx59 = multm_reduce_mulsc_mulb_yoc59 & multm_reduce_mulsc_mulb_ps59;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx60 = multm_reduce_mulsc_mulb_yoc60 & multm_reduce_mulsc_mulb_ps60;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx61 = multm_reduce_mulsc_mulb_yoc61 & multm_reduce_mulsc_mulb_ps61;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx62 = multm_reduce_mulsc_mulb_yoc62 & multm_reduce_mulsc_mulb_ps62;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx63 = multm_reduce_mulsc_mulb_yoc63 & multm_reduce_mulsc_mulb_ps63;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx64 = multm_reduce_mulsc_mulb_yoc64 & multm_reduce_mulsc_mulb_ps64;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx65 = multm_reduce_mulsc_mulb_yoc65 & multm_reduce_mulsc_mulb_ps65;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx66 = multm_reduce_mulsc_mulb_yoc66 & multm_reduce_mulsc_mulb_ps66;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx67 = multm_reduce_mulsc_mulb_yoc67 & multm_reduce_mulsc_mulb_ps67;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx68 = multm_reduce_mulsc_mulb_yoc68 & multm_reduce_mulsc_mulb_ps68;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx69 = multm_reduce_mulsc_mulb_yoc69 & multm_reduce_mulsc_mulb_ps69;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx70 = multm_reduce_mulsc_mulb_yoc70 & multm_reduce_mulsc_mulb_ps70;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx71 = multm_reduce_mulsc_mulb_yoc71 & multm_reduce_mulsc_mulb_ps71;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx72 = multm_reduce_mulsc_mulb_yoc72 & multm_reduce_mulsc_mulb_ps72;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx73 = multm_reduce_mulsc_mulb_yoc73 & multm_reduce_mulsc_mulb_ps73;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx74 = multm_reduce_mulsc_mulb_yoc74 & multm_reduce_mulsc_mulb_ps74;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx75 = multm_reduce_mulsc_mulb_yoc75 & multm_reduce_mulsc_mulb_ps75;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx76 = multm_reduce_mulsc_mulb_yoc76 & multm_reduce_mulsc_mulb_ps76;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx77 = multm_reduce_mulsc_mulb_yoc77 & multm_reduce_mulsc_mulb_ps77;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx78 = multm_reduce_mulsc_mulb_yoc78 & multm_reduce_mulsc_mulb_ps78;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx79 = multm_reduce_mulsc_mulb_yoc79 & multm_reduce_mulsc_mulb_ps79;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx80 = multm_reduce_mulsc_mulb_yoc80 & multm_reduce_mulsc_mulb_ps80;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx81 = multm_reduce_mulsc_mulb_yoc81 & multm_reduce_mulsc_mulb_ps81;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx82 = multm_reduce_mulsc_mulb_yoc82 & multm_reduce_mulsc_mulb_ps82;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx83 = multm_reduce_mulsc_mulb_yoc83 & multm_reduce_mulsc_mulb_ps83;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx84 = multm_reduce_mulsc_mulb_yoc84 & multm_reduce_mulsc_mulb_ps84;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx85 = multm_reduce_mulsc_mulb_yoc85 & multm_reduce_mulsc_mulb_ps85;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx86 = multm_reduce_mulsc_mulb_yoc86 & multm_reduce_mulsc_mulb_ps86;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx87 = multm_reduce_mulsc_mulb_yoc87 & multm_reduce_mulsc_mulb_ps87;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx88 = multm_reduce_mulsc_mulb_yoc88 & multm_reduce_mulsc_mulb_ps88;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx89 = multm_reduce_mulsc_mulb_yoc89 & multm_reduce_mulsc_mulb_ps89;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx90 = multm_reduce_mulsc_mulb_yoc90 & multm_reduce_mulsc_mulb_ps90;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx91 = multm_reduce_mulsc_mulb_yoc91 & multm_reduce_mulsc_mulb_ps91;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx92 = multm_reduce_mulsc_mulb_yoc92 & multm_reduce_mulsc_mulb_ps92;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx93 = multm_reduce_mulsc_mulb_yoc93 & multm_reduce_mulsc_mulb_ps93;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx94 = multm_reduce_mulsc_mulb_yoc94 & multm_reduce_mulsc_mulb_ps94;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx95 = multm_reduce_mulsc_mulb_yoc95 & multm_reduce_mulsc_mulb_ps95;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx96 = multm_reduce_mulsc_mulb_yoc96 & multm_reduce_mulsc_mulb_ps96;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx97 = multm_reduce_mulsc_mulb_yoc97 & multm_reduce_mulsc_mulb_ps97;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx98 = multm_reduce_mulsc_mulb_yoc98 & multm_reduce_mulsc_mulb_ps98;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx99 = multm_reduce_mulsc_mulb_yoc99 & multm_reduce_mulsc_mulb_ps99;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx100 = multm_reduce_mulsc_mulb_yoc100 & multm_reduce_mulsc_mulb_ps100;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx101 = multm_reduce_mulsc_mulb_yoc101 & multm_reduce_mulsc_mulb_ps101;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx102 = multm_reduce_mulsc_mulb_yoc102 & multm_reduce_mulsc_mulb_ps102;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx103 = multm_reduce_mulsc_mulb_yoc103 & multm_reduce_mulsc_mulb_ps103;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx104 = multm_reduce_mulsc_mulb_yoc104 & multm_reduce_mulsc_mulb_ps104;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx105 = multm_reduce_mulsc_mulb_yoc105 & multm_reduce_mulsc_mulb_ps105;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx106 = multm_reduce_mulsc_mulb_yoc106 & multm_reduce_mulsc_mulb_ps106;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx107 = multm_reduce_mulsc_mulb_yoc107 & multm_reduce_mulsc_mulb_ps107;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx108 = multm_reduce_mulsc_mulb_yoc108 & multm_reduce_mulsc_mulb_ps108;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx109 = multm_reduce_mulsc_mulb_yoc109 & multm_reduce_mulsc_mulb_ps109;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx110 = multm_reduce_mulsc_mulb_yoc110 & multm_reduce_mulsc_mulb_ps110;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx111 = multm_reduce_mulsc_mulb_yoc111 & multm_reduce_mulsc_mulb_ps111;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx112 = multm_reduce_mulsc_mulb_yoc112 & multm_reduce_mulsc_mulb_ps112;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx113 = multm_reduce_mulsc_mulb_yoc113 & multm_reduce_mulsc_mulb_ps113;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx114 = multm_reduce_mulsc_mulb_yoc114 & multm_reduce_mulsc_mulb_ps114;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx115 = multm_reduce_mulsc_mulb_yoc115 & multm_reduce_mulsc_mulb_ps115;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx116 = multm_reduce_mulsc_mulb_yoc116 & multm_reduce_mulsc_mulb_ps116;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx117 = multm_reduce_mulsc_mulb_yoc117 & multm_reduce_mulsc_mulb_ps117;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx118 = multm_reduce_mulsc_mulb_yoc118 & multm_reduce_mulsc_mulb_ps118;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx119 = multm_reduce_mulsc_mulb_yoc119 & multm_reduce_mulsc_mulb_ps119;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx120 = multm_reduce_mulsc_mulb_yoc120 & multm_reduce_mulsc_mulb_ps120;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx121 = multm_reduce_mulsc_mulb_yoc121 & multm_reduce_mulsc_mulb_ps121;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx122 = multm_reduce_mulsc_mulb_yoc122 & multm_reduce_mulsc_mulb_ps122;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx123 = multm_reduce_mulsc_mulb_yoc123 & multm_reduce_mulsc_mulb_ps123;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx124 = multm_reduce_mulsc_mulb_yoc124 & multm_reduce_mulsc_mulb_ps124;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx125 = multm_reduce_mulsc_mulb_yoc125 & multm_reduce_mulsc_mulb_ps125;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx126 = multm_reduce_mulsc_mulb_yoc126 & multm_reduce_mulsc_mulb_ps126;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx127 = multm_reduce_mulsc_mulb_yoc127 & multm_reduce_mulsc_mulb_ps127;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx128 = multm_reduce_mulsc_mulb_yoc128 & multm_reduce_mulsc_mulb_ps128;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx129 = multm_reduce_mulsc_mulb_yoc129 & multm_reduce_mulsc_mulb_ps129;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx130 = multm_reduce_mulsc_mulb_yoc130 & multm_reduce_mulsc_mulb_ps130;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx131 = multm_reduce_mulsc_mulb_yoc131 & multm_reduce_mulsc_mulb_ps131;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx132 = multm_reduce_mulsc_mulb_yoc132 & multm_reduce_mulsc_mulb_ps132;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx133 = multm_reduce_mulsc_mulb_yoc133 & multm_reduce_mulsc_mulb_ps133;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx134 = multm_reduce_mulsc_mulb_yoc134 & multm_reduce_mulsc_mulb_ps134;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx135 = multm_reduce_mulsc_mulb_yoc135 & multm_reduce_mulsc_mulb_ps135;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx136 = multm_reduce_mulsc_mulb_yoc136 & multm_reduce_mulsc_mulb_ps136;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx137 = multm_reduce_mulsc_mulb_yoc137 & multm_reduce_mulsc_mulb_ps137;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx138 = multm_reduce_mulsc_mulb_yoc138 & multm_reduce_mulsc_mulb_ps138;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx139 = multm_reduce_mulsc_mulb_yoc139 & multm_reduce_mulsc_mulb_ps139;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx140 = multm_reduce_mulsc_mulb_yoc140 & multm_reduce_mulsc_mulb_ps140;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx141 = multm_reduce_mulsc_mulb_yoc141 & multm_reduce_mulsc_mulb_ps141;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx142 = multm_reduce_mulsc_mulb_yoc142 & multm_reduce_mulsc_mulb_ps142;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx143 = multm_reduce_mulsc_mulb_yoc143 & multm_reduce_mulsc_mulb_ps143;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx144 = multm_reduce_mulsc_mulb_yoc144 & multm_reduce_mulsc_mulb_ps144;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx145 = multm_reduce_mulsc_mulb_yoc145 & multm_reduce_mulsc_mulb_ps145;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx146 = multm_reduce_mulsc_mulb_yoc146 & multm_reduce_mulsc_mulb_ps146;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx147 = multm_reduce_mulsc_mulb_yoc147 & multm_reduce_mulsc_mulb_ps147;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx148 = multm_reduce_mulsc_mulb_yoc148 & multm_reduce_mulsc_mulb_ps148;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx149 = multm_reduce_mulsc_mulb_yoc149 & multm_reduce_mulsc_mulb_ps149;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx150 = multm_reduce_mulsc_mulb_yoc150 & multm_reduce_mulsc_mulb_ps150;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx151 = multm_reduce_mulsc_mulb_yoc151 & multm_reduce_mulsc_mulb_ps151;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx152 = multm_reduce_mulsc_mulb_yoc152 & multm_reduce_mulsc_mulb_ps152;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx153 = multm_reduce_mulsc_mulb_yoc153 & multm_reduce_mulsc_mulb_ps153;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx154 = multm_reduce_mulsc_mulb_yoc154 & multm_reduce_mulsc_mulb_ps154;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx155 = multm_reduce_mulsc_mulb_yoc155 & multm_reduce_mulsc_mulb_ps155;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx156 = multm_reduce_mulsc_mulb_yoc156 & multm_reduce_mulsc_mulb_ps156;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx157 = multm_reduce_mulsc_mulb_yoc157 & multm_reduce_mulsc_mulb_ps157;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx158 = multm_reduce_mulsc_mulb_yoc158 & multm_reduce_mulsc_mulb_ps158;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx159 = multm_reduce_mulsc_mulb_yoc159 & multm_reduce_mulsc_mulb_ps159;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx160 = multm_reduce_mulsc_mulb_yoc160 & multm_reduce_mulsc_mulb_ps160;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx161 = multm_reduce_mulsc_mulb_yoc161 & multm_reduce_mulsc_mulb_ps161;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx162 = multm_reduce_mulsc_mulb_yoc162 & multm_reduce_mulsc_mulb_ps162;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx163 = multm_reduce_mulsc_mulb_yoc163 & multm_reduce_mulsc_mulb_ps163;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx164 = multm_reduce_mulsc_mulb_yoc164 & multm_reduce_mulsc_mulb_ps164;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx165 = multm_reduce_mulsc_mulb_yoc165 & multm_reduce_mulsc_mulb_ps165;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx166 = multm_reduce_mulsc_mulb_yoc166 & multm_reduce_mulsc_mulb_ps166;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx167 = multm_reduce_mulsc_mulb_yoc167 & multm_reduce_mulsc_mulb_ps167;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx168 = multm_reduce_mulsc_mulb_yoc168 & multm_reduce_mulsc_mulb_ps168;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx169 = multm_reduce_mulsc_mulb_yoc169 & multm_reduce_mulsc_mulb_ps169;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx170 = multm_reduce_mulsc_mulb_yoc170 & multm_reduce_mulsc_mulb_ps170;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx171 = multm_reduce_mulsc_mulb_yoc171 & multm_reduce_mulsc_mulb_ps171;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx172 = multm_reduce_mulsc_mulb_yoc172 & multm_reduce_mulsc_mulb_ps172;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx173 = multm_reduce_mulsc_mulb_yoc173 & multm_reduce_mulsc_mulb_ps173;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx174 = multm_reduce_mulsc_mulb_yoc174 & multm_reduce_mulsc_mulb_ps174;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx175 = multm_reduce_mulsc_mulb_yoc175 & multm_reduce_mulsc_mulb_ps175;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx176 = multm_reduce_mulsc_mulb_yoc176 & multm_reduce_mulsc_mulb_ps176;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx177 = multm_reduce_mulsc_mulb_yoc177 & multm_reduce_mulsc_mulb_ps177;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx178 = multm_reduce_mulsc_mulb_yoc178 & multm_reduce_mulsc_mulb_ps178;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx179 = multm_reduce_mulsc_mulb_yoc179 & multm_reduce_mulsc_mulb_ps179;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx180 = multm_reduce_mulsc_mulb_yoc180 & multm_reduce_mulsc_mulb_ps180;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx181 = multm_reduce_mulsc_mulb_yoc181 & multm_reduce_mulsc_mulb_ps181;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wx182 = multm_reduce_mulsc_mulb_yoc182 & multm_reduce_mulsc_mulb_ps182;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy0 = multm_reduce_mulsc_mulb_yoc0 & multm_reduce_mulsc_mulb_pc0;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy1 = multm_reduce_mulsc_mulb_yoc1 & multm_reduce_mulsc_mulb_pc1;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy2 = multm_reduce_mulsc_mulb_yoc2 & multm_reduce_mulsc_mulb_pc2;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy3 = multm_reduce_mulsc_mulb_yoc3 & multm_reduce_mulsc_mulb_pc3;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy4 = multm_reduce_mulsc_mulb_yoc4 & multm_reduce_mulsc_mulb_pc4;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy5 = multm_reduce_mulsc_mulb_yoc5 & multm_reduce_mulsc_mulb_pc5;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy6 = multm_reduce_mulsc_mulb_yoc6 & multm_reduce_mulsc_mulb_pc6;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy7 = multm_reduce_mulsc_mulb_yoc7 & multm_reduce_mulsc_mulb_pc7;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy8 = multm_reduce_mulsc_mulb_yoc8 & multm_reduce_mulsc_mulb_pc8;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy9 = multm_reduce_mulsc_mulb_yoc9 & multm_reduce_mulsc_mulb_pc9;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy10 = multm_reduce_mulsc_mulb_yoc10 & multm_reduce_mulsc_mulb_pc10;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy11 = multm_reduce_mulsc_mulb_yoc11 & multm_reduce_mulsc_mulb_pc11;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy12 = multm_reduce_mulsc_mulb_yoc12 & multm_reduce_mulsc_mulb_pc12;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy13 = multm_reduce_mulsc_mulb_yoc13 & multm_reduce_mulsc_mulb_pc13;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy14 = multm_reduce_mulsc_mulb_yoc14 & multm_reduce_mulsc_mulb_pc14;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy15 = multm_reduce_mulsc_mulb_yoc15 & multm_reduce_mulsc_mulb_pc15;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy16 = multm_reduce_mulsc_mulb_yoc16 & multm_reduce_mulsc_mulb_pc16;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy17 = multm_reduce_mulsc_mulb_yoc17 & multm_reduce_mulsc_mulb_pc17;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy18 = multm_reduce_mulsc_mulb_yoc18 & multm_reduce_mulsc_mulb_pc18;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy19 = multm_reduce_mulsc_mulb_yoc19 & multm_reduce_mulsc_mulb_pc19;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy20 = multm_reduce_mulsc_mulb_yoc20 & multm_reduce_mulsc_mulb_pc20;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy21 = multm_reduce_mulsc_mulb_yoc21 & multm_reduce_mulsc_mulb_pc21;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy22 = multm_reduce_mulsc_mulb_yoc22 & multm_reduce_mulsc_mulb_pc22;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy23 = multm_reduce_mulsc_mulb_yoc23 & multm_reduce_mulsc_mulb_pc23;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy24 = multm_reduce_mulsc_mulb_yoc24 & multm_reduce_mulsc_mulb_pc24;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy25 = multm_reduce_mulsc_mulb_yoc25 & multm_reduce_mulsc_mulb_pc25;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy26 = multm_reduce_mulsc_mulb_yoc26 & multm_reduce_mulsc_mulb_pc26;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy27 = multm_reduce_mulsc_mulb_yoc27 & multm_reduce_mulsc_mulb_pc27;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy28 = multm_reduce_mulsc_mulb_yoc28 & multm_reduce_mulsc_mulb_pc28;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy29 = multm_reduce_mulsc_mulb_yoc29 & multm_reduce_mulsc_mulb_pc29;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy30 = multm_reduce_mulsc_mulb_yoc30 & multm_reduce_mulsc_mulb_pc30;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy31 = multm_reduce_mulsc_mulb_yoc31 & multm_reduce_mulsc_mulb_pc31;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy32 = multm_reduce_mulsc_mulb_yoc32 & multm_reduce_mulsc_mulb_pc32;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy33 = multm_reduce_mulsc_mulb_yoc33 & multm_reduce_mulsc_mulb_pc33;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy34 = multm_reduce_mulsc_mulb_yoc34 & multm_reduce_mulsc_mulb_pc34;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy35 = multm_reduce_mulsc_mulb_yoc35 & multm_reduce_mulsc_mulb_pc35;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy36 = multm_reduce_mulsc_mulb_yoc36 & multm_reduce_mulsc_mulb_pc36;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy37 = multm_reduce_mulsc_mulb_yoc37 & multm_reduce_mulsc_mulb_pc37;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy38 = multm_reduce_mulsc_mulb_yoc38 & multm_reduce_mulsc_mulb_pc38;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy39 = multm_reduce_mulsc_mulb_yoc39 & multm_reduce_mulsc_mulb_pc39;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy40 = multm_reduce_mulsc_mulb_yoc40 & multm_reduce_mulsc_mulb_pc40;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy41 = multm_reduce_mulsc_mulb_yoc41 & multm_reduce_mulsc_mulb_pc41;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy42 = multm_reduce_mulsc_mulb_yoc42 & multm_reduce_mulsc_mulb_pc42;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy43 = multm_reduce_mulsc_mulb_yoc43 & multm_reduce_mulsc_mulb_pc43;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy44 = multm_reduce_mulsc_mulb_yoc44 & multm_reduce_mulsc_mulb_pc44;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy45 = multm_reduce_mulsc_mulb_yoc45 & multm_reduce_mulsc_mulb_pc45;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy46 = multm_reduce_mulsc_mulb_yoc46 & multm_reduce_mulsc_mulb_pc46;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy47 = multm_reduce_mulsc_mulb_yoc47 & multm_reduce_mulsc_mulb_pc47;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy48 = multm_reduce_mulsc_mulb_yoc48 & multm_reduce_mulsc_mulb_pc48;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy49 = multm_reduce_mulsc_mulb_yoc49 & multm_reduce_mulsc_mulb_pc49;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy50 = multm_reduce_mulsc_mulb_yoc50 & multm_reduce_mulsc_mulb_pc50;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy51 = multm_reduce_mulsc_mulb_yoc51 & multm_reduce_mulsc_mulb_pc51;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy52 = multm_reduce_mulsc_mulb_yoc52 & multm_reduce_mulsc_mulb_pc52;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy53 = multm_reduce_mulsc_mulb_yoc53 & multm_reduce_mulsc_mulb_pc53;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy54 = multm_reduce_mulsc_mulb_yoc54 & multm_reduce_mulsc_mulb_pc54;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy55 = multm_reduce_mulsc_mulb_yoc55 & multm_reduce_mulsc_mulb_pc55;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy56 = multm_reduce_mulsc_mulb_yoc56 & multm_reduce_mulsc_mulb_pc56;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy57 = multm_reduce_mulsc_mulb_yoc57 & multm_reduce_mulsc_mulb_pc57;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy58 = multm_reduce_mulsc_mulb_yoc58 & multm_reduce_mulsc_mulb_pc58;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy59 = multm_reduce_mulsc_mulb_yoc59 & multm_reduce_mulsc_mulb_pc59;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy60 = multm_reduce_mulsc_mulb_yoc60 & multm_reduce_mulsc_mulb_pc60;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy61 = multm_reduce_mulsc_mulb_yoc61 & multm_reduce_mulsc_mulb_pc61;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy62 = multm_reduce_mulsc_mulb_yoc62 & multm_reduce_mulsc_mulb_pc62;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy63 = multm_reduce_mulsc_mulb_yoc63 & multm_reduce_mulsc_mulb_pc63;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy64 = multm_reduce_mulsc_mulb_yoc64 & multm_reduce_mulsc_mulb_pc64;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy65 = multm_reduce_mulsc_mulb_yoc65 & multm_reduce_mulsc_mulb_pc65;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy66 = multm_reduce_mulsc_mulb_yoc66 & multm_reduce_mulsc_mulb_pc66;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy67 = multm_reduce_mulsc_mulb_yoc67 & multm_reduce_mulsc_mulb_pc67;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy68 = multm_reduce_mulsc_mulb_yoc68 & multm_reduce_mulsc_mulb_pc68;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy69 = multm_reduce_mulsc_mulb_yoc69 & multm_reduce_mulsc_mulb_pc69;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy70 = multm_reduce_mulsc_mulb_yoc70 & multm_reduce_mulsc_mulb_pc70;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy71 = multm_reduce_mulsc_mulb_yoc71 & multm_reduce_mulsc_mulb_pc71;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy72 = multm_reduce_mulsc_mulb_yoc72 & multm_reduce_mulsc_mulb_pc72;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy73 = multm_reduce_mulsc_mulb_yoc73 & multm_reduce_mulsc_mulb_pc73;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy74 = multm_reduce_mulsc_mulb_yoc74 & multm_reduce_mulsc_mulb_pc74;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy75 = multm_reduce_mulsc_mulb_yoc75 & multm_reduce_mulsc_mulb_pc75;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy76 = multm_reduce_mulsc_mulb_yoc76 & multm_reduce_mulsc_mulb_pc76;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy77 = multm_reduce_mulsc_mulb_yoc77 & multm_reduce_mulsc_mulb_pc77;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy78 = multm_reduce_mulsc_mulb_yoc78 & multm_reduce_mulsc_mulb_pc78;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy79 = multm_reduce_mulsc_mulb_yoc79 & multm_reduce_mulsc_mulb_pc79;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy80 = multm_reduce_mulsc_mulb_yoc80 & multm_reduce_mulsc_mulb_pc80;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy81 = multm_reduce_mulsc_mulb_yoc81 & multm_reduce_mulsc_mulb_pc81;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy82 = multm_reduce_mulsc_mulb_yoc82 & multm_reduce_mulsc_mulb_pc82;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy83 = multm_reduce_mulsc_mulb_yoc83 & multm_reduce_mulsc_mulb_pc83;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy84 = multm_reduce_mulsc_mulb_yoc84 & multm_reduce_mulsc_mulb_pc84;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy85 = multm_reduce_mulsc_mulb_yoc85 & multm_reduce_mulsc_mulb_pc85;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy86 = multm_reduce_mulsc_mulb_yoc86 & multm_reduce_mulsc_mulb_pc86;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy87 = multm_reduce_mulsc_mulb_yoc87 & multm_reduce_mulsc_mulb_pc87;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy88 = multm_reduce_mulsc_mulb_yoc88 & multm_reduce_mulsc_mulb_pc88;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy89 = multm_reduce_mulsc_mulb_yoc89 & multm_reduce_mulsc_mulb_pc89;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy90 = multm_reduce_mulsc_mulb_yoc90 & multm_reduce_mulsc_mulb_pc90;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy91 = multm_reduce_mulsc_mulb_yoc91 & multm_reduce_mulsc_mulb_pc91;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy92 = multm_reduce_mulsc_mulb_yoc92 & multm_reduce_mulsc_mulb_pc92;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy93 = multm_reduce_mulsc_mulb_yoc93 & multm_reduce_mulsc_mulb_pc93;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy94 = multm_reduce_mulsc_mulb_yoc94 & multm_reduce_mulsc_mulb_pc94;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy95 = multm_reduce_mulsc_mulb_yoc95 & multm_reduce_mulsc_mulb_pc95;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy96 = multm_reduce_mulsc_mulb_yoc96 & multm_reduce_mulsc_mulb_pc96;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy97 = multm_reduce_mulsc_mulb_yoc97 & multm_reduce_mulsc_mulb_pc97;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy98 = multm_reduce_mulsc_mulb_yoc98 & multm_reduce_mulsc_mulb_pc98;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy99 = multm_reduce_mulsc_mulb_yoc99 & multm_reduce_mulsc_mulb_pc99;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy100 = multm_reduce_mulsc_mulb_yoc100 & multm_reduce_mulsc_mulb_pc100;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy101 = multm_reduce_mulsc_mulb_yoc101 & multm_reduce_mulsc_mulb_pc101;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy102 = multm_reduce_mulsc_mulb_yoc102 & multm_reduce_mulsc_mulb_pc102;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy103 = multm_reduce_mulsc_mulb_yoc103 & multm_reduce_mulsc_mulb_pc103;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy104 = multm_reduce_mulsc_mulb_yoc104 & multm_reduce_mulsc_mulb_pc104;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy105 = multm_reduce_mulsc_mulb_yoc105 & multm_reduce_mulsc_mulb_pc105;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy106 = multm_reduce_mulsc_mulb_yoc106 & multm_reduce_mulsc_mulb_pc106;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy107 = multm_reduce_mulsc_mulb_yoc107 & multm_reduce_mulsc_mulb_pc107;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy108 = multm_reduce_mulsc_mulb_yoc108 & multm_reduce_mulsc_mulb_pc108;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy109 = multm_reduce_mulsc_mulb_yoc109 & multm_reduce_mulsc_mulb_pc109;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy110 = multm_reduce_mulsc_mulb_yoc110 & multm_reduce_mulsc_mulb_pc110;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy111 = multm_reduce_mulsc_mulb_yoc111 & multm_reduce_mulsc_mulb_pc111;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy112 = multm_reduce_mulsc_mulb_yoc112 & multm_reduce_mulsc_mulb_pc112;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy113 = multm_reduce_mulsc_mulb_yoc113 & multm_reduce_mulsc_mulb_pc113;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy114 = multm_reduce_mulsc_mulb_yoc114 & multm_reduce_mulsc_mulb_pc114;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy115 = multm_reduce_mulsc_mulb_yoc115 & multm_reduce_mulsc_mulb_pc115;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy116 = multm_reduce_mulsc_mulb_yoc116 & multm_reduce_mulsc_mulb_pc116;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy117 = multm_reduce_mulsc_mulb_yoc117 & multm_reduce_mulsc_mulb_pc117;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy118 = multm_reduce_mulsc_mulb_yoc118 & multm_reduce_mulsc_mulb_pc118;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy119 = multm_reduce_mulsc_mulb_yoc119 & multm_reduce_mulsc_mulb_pc119;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy120 = multm_reduce_mulsc_mulb_yoc120 & multm_reduce_mulsc_mulb_pc120;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy121 = multm_reduce_mulsc_mulb_yoc121 & multm_reduce_mulsc_mulb_pc121;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy122 = multm_reduce_mulsc_mulb_yoc122 & multm_reduce_mulsc_mulb_pc122;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy123 = multm_reduce_mulsc_mulb_yoc123 & multm_reduce_mulsc_mulb_pc123;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy124 = multm_reduce_mulsc_mulb_yoc124 & multm_reduce_mulsc_mulb_pc124;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy125 = multm_reduce_mulsc_mulb_yoc125 & multm_reduce_mulsc_mulb_pc125;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy126 = multm_reduce_mulsc_mulb_yoc126 & multm_reduce_mulsc_mulb_pc126;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy127 = multm_reduce_mulsc_mulb_yoc127 & multm_reduce_mulsc_mulb_pc127;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy128 = multm_reduce_mulsc_mulb_yoc128 & multm_reduce_mulsc_mulb_pc128;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy129 = multm_reduce_mulsc_mulb_yoc129 & multm_reduce_mulsc_mulb_pc129;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy130 = multm_reduce_mulsc_mulb_yoc130 & multm_reduce_mulsc_mulb_pc130;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy131 = multm_reduce_mulsc_mulb_yoc131 & multm_reduce_mulsc_mulb_pc131;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy132 = multm_reduce_mulsc_mulb_yoc132 & multm_reduce_mulsc_mulb_pc132;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy133 = multm_reduce_mulsc_mulb_yoc133 & multm_reduce_mulsc_mulb_pc133;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy134 = multm_reduce_mulsc_mulb_yoc134 & multm_reduce_mulsc_mulb_pc134;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy135 = multm_reduce_mulsc_mulb_yoc135 & multm_reduce_mulsc_mulb_pc135;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy136 = multm_reduce_mulsc_mulb_yoc136 & multm_reduce_mulsc_mulb_pc136;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy137 = multm_reduce_mulsc_mulb_yoc137 & multm_reduce_mulsc_mulb_pc137;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy138 = multm_reduce_mulsc_mulb_yoc138 & multm_reduce_mulsc_mulb_pc138;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy139 = multm_reduce_mulsc_mulb_yoc139 & multm_reduce_mulsc_mulb_pc139;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy140 = multm_reduce_mulsc_mulb_yoc140 & multm_reduce_mulsc_mulb_pc140;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy141 = multm_reduce_mulsc_mulb_yoc141 & multm_reduce_mulsc_mulb_pc141;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy142 = multm_reduce_mulsc_mulb_yoc142 & multm_reduce_mulsc_mulb_pc142;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy143 = multm_reduce_mulsc_mulb_yoc143 & multm_reduce_mulsc_mulb_pc143;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy144 = multm_reduce_mulsc_mulb_yoc144 & multm_reduce_mulsc_mulb_pc144;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy145 = multm_reduce_mulsc_mulb_yoc145 & multm_reduce_mulsc_mulb_pc145;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy146 = multm_reduce_mulsc_mulb_yoc146 & multm_reduce_mulsc_mulb_pc146;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy147 = multm_reduce_mulsc_mulb_yoc147 & multm_reduce_mulsc_mulb_pc147;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy148 = multm_reduce_mulsc_mulb_yoc148 & multm_reduce_mulsc_mulb_pc148;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy149 = multm_reduce_mulsc_mulb_yoc149 & multm_reduce_mulsc_mulb_pc149;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy150 = multm_reduce_mulsc_mulb_yoc150 & multm_reduce_mulsc_mulb_pc150;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy151 = multm_reduce_mulsc_mulb_yoc151 & multm_reduce_mulsc_mulb_pc151;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy152 = multm_reduce_mulsc_mulb_yoc152 & multm_reduce_mulsc_mulb_pc152;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy153 = multm_reduce_mulsc_mulb_yoc153 & multm_reduce_mulsc_mulb_pc153;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy154 = multm_reduce_mulsc_mulb_yoc154 & multm_reduce_mulsc_mulb_pc154;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy155 = multm_reduce_mulsc_mulb_yoc155 & multm_reduce_mulsc_mulb_pc155;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy156 = multm_reduce_mulsc_mulb_yoc156 & multm_reduce_mulsc_mulb_pc156;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy157 = multm_reduce_mulsc_mulb_yoc157 & multm_reduce_mulsc_mulb_pc157;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy158 = multm_reduce_mulsc_mulb_yoc158 & multm_reduce_mulsc_mulb_pc158;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy159 = multm_reduce_mulsc_mulb_yoc159 & multm_reduce_mulsc_mulb_pc159;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy160 = multm_reduce_mulsc_mulb_yoc160 & multm_reduce_mulsc_mulb_pc160;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy161 = multm_reduce_mulsc_mulb_yoc161 & multm_reduce_mulsc_mulb_pc161;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy162 = multm_reduce_mulsc_mulb_yoc162 & multm_reduce_mulsc_mulb_pc162;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy163 = multm_reduce_mulsc_mulb_yoc163 & multm_reduce_mulsc_mulb_pc163;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy164 = multm_reduce_mulsc_mulb_yoc164 & multm_reduce_mulsc_mulb_pc164;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy165 = multm_reduce_mulsc_mulb_yoc165 & multm_reduce_mulsc_mulb_pc165;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy166 = multm_reduce_mulsc_mulb_yoc166 & multm_reduce_mulsc_mulb_pc166;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy167 = multm_reduce_mulsc_mulb_yoc167 & multm_reduce_mulsc_mulb_pc167;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy168 = multm_reduce_mulsc_mulb_yoc168 & multm_reduce_mulsc_mulb_pc168;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy169 = multm_reduce_mulsc_mulb_yoc169 & multm_reduce_mulsc_mulb_pc169;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy170 = multm_reduce_mulsc_mulb_yoc170 & multm_reduce_mulsc_mulb_pc170;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy171 = multm_reduce_mulsc_mulb_yoc171 & multm_reduce_mulsc_mulb_pc171;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy172 = multm_reduce_mulsc_mulb_yoc172 & multm_reduce_mulsc_mulb_pc172;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy173 = multm_reduce_mulsc_mulb_yoc173 & multm_reduce_mulsc_mulb_pc173;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy174 = multm_reduce_mulsc_mulb_yoc174 & multm_reduce_mulsc_mulb_pc174;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy175 = multm_reduce_mulsc_mulb_yoc175 & multm_reduce_mulsc_mulb_pc175;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy176 = multm_reduce_mulsc_mulb_yoc176 & multm_reduce_mulsc_mulb_pc176;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy177 = multm_reduce_mulsc_mulb_yoc177 & multm_reduce_mulsc_mulb_pc177;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy178 = multm_reduce_mulsc_mulb_yoc178 & multm_reduce_mulsc_mulb_pc178;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy179 = multm_reduce_mulsc_mulb_yoc179 & multm_reduce_mulsc_mulb_pc179;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy180 = multm_reduce_mulsc_mulb_yoc180 & multm_reduce_mulsc_mulb_pc180;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy181 = multm_reduce_mulsc_mulb_yoc181 & multm_reduce_mulsc_mulb_pc181;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_wy182 = multm_reduce_mulsc_mulb_yoc182 & multm_reduce_mulsc_mulb_pc182;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy0 = multm_reduce_mulsc_mulb_ps0 & multm_reduce_mulsc_mulb_pc0;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy1 = multm_reduce_mulsc_mulb_ps1 & multm_reduce_mulsc_mulb_pc1;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy2 = multm_reduce_mulsc_mulb_ps2 & multm_reduce_mulsc_mulb_pc2;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy3 = multm_reduce_mulsc_mulb_ps3 & multm_reduce_mulsc_mulb_pc3;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy4 = multm_reduce_mulsc_mulb_ps4 & multm_reduce_mulsc_mulb_pc4;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy5 = multm_reduce_mulsc_mulb_ps5 & multm_reduce_mulsc_mulb_pc5;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy6 = multm_reduce_mulsc_mulb_ps6 & multm_reduce_mulsc_mulb_pc6;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy7 = multm_reduce_mulsc_mulb_ps7 & multm_reduce_mulsc_mulb_pc7;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy8 = multm_reduce_mulsc_mulb_ps8 & multm_reduce_mulsc_mulb_pc8;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy9 = multm_reduce_mulsc_mulb_ps9 & multm_reduce_mulsc_mulb_pc9;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy10 = multm_reduce_mulsc_mulb_ps10 & multm_reduce_mulsc_mulb_pc10;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy11 = multm_reduce_mulsc_mulb_ps11 & multm_reduce_mulsc_mulb_pc11;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy12 = multm_reduce_mulsc_mulb_ps12 & multm_reduce_mulsc_mulb_pc12;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy13 = multm_reduce_mulsc_mulb_ps13 & multm_reduce_mulsc_mulb_pc13;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy14 = multm_reduce_mulsc_mulb_ps14 & multm_reduce_mulsc_mulb_pc14;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy15 = multm_reduce_mulsc_mulb_ps15 & multm_reduce_mulsc_mulb_pc15;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy16 = multm_reduce_mulsc_mulb_ps16 & multm_reduce_mulsc_mulb_pc16;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy17 = multm_reduce_mulsc_mulb_ps17 & multm_reduce_mulsc_mulb_pc17;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy18 = multm_reduce_mulsc_mulb_ps18 & multm_reduce_mulsc_mulb_pc18;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy19 = multm_reduce_mulsc_mulb_ps19 & multm_reduce_mulsc_mulb_pc19;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy20 = multm_reduce_mulsc_mulb_ps20 & multm_reduce_mulsc_mulb_pc20;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy21 = multm_reduce_mulsc_mulb_ps21 & multm_reduce_mulsc_mulb_pc21;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy22 = multm_reduce_mulsc_mulb_ps22 & multm_reduce_mulsc_mulb_pc22;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy23 = multm_reduce_mulsc_mulb_ps23 & multm_reduce_mulsc_mulb_pc23;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy24 = multm_reduce_mulsc_mulb_ps24 & multm_reduce_mulsc_mulb_pc24;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy25 = multm_reduce_mulsc_mulb_ps25 & multm_reduce_mulsc_mulb_pc25;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy26 = multm_reduce_mulsc_mulb_ps26 & multm_reduce_mulsc_mulb_pc26;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy27 = multm_reduce_mulsc_mulb_ps27 & multm_reduce_mulsc_mulb_pc27;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy28 = multm_reduce_mulsc_mulb_ps28 & multm_reduce_mulsc_mulb_pc28;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy29 = multm_reduce_mulsc_mulb_ps29 & multm_reduce_mulsc_mulb_pc29;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy30 = multm_reduce_mulsc_mulb_ps30 & multm_reduce_mulsc_mulb_pc30;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy31 = multm_reduce_mulsc_mulb_ps31 & multm_reduce_mulsc_mulb_pc31;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy32 = multm_reduce_mulsc_mulb_ps32 & multm_reduce_mulsc_mulb_pc32;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy33 = multm_reduce_mulsc_mulb_ps33 & multm_reduce_mulsc_mulb_pc33;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy34 = multm_reduce_mulsc_mulb_ps34 & multm_reduce_mulsc_mulb_pc34;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy35 = multm_reduce_mulsc_mulb_ps35 & multm_reduce_mulsc_mulb_pc35;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy36 = multm_reduce_mulsc_mulb_ps36 & multm_reduce_mulsc_mulb_pc36;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy37 = multm_reduce_mulsc_mulb_ps37 & multm_reduce_mulsc_mulb_pc37;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy38 = multm_reduce_mulsc_mulb_ps38 & multm_reduce_mulsc_mulb_pc38;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy39 = multm_reduce_mulsc_mulb_ps39 & multm_reduce_mulsc_mulb_pc39;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy40 = multm_reduce_mulsc_mulb_ps40 & multm_reduce_mulsc_mulb_pc40;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy41 = multm_reduce_mulsc_mulb_ps41 & multm_reduce_mulsc_mulb_pc41;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy42 = multm_reduce_mulsc_mulb_ps42 & multm_reduce_mulsc_mulb_pc42;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy43 = multm_reduce_mulsc_mulb_ps43 & multm_reduce_mulsc_mulb_pc43;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy44 = multm_reduce_mulsc_mulb_ps44 & multm_reduce_mulsc_mulb_pc44;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy45 = multm_reduce_mulsc_mulb_ps45 & multm_reduce_mulsc_mulb_pc45;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy46 = multm_reduce_mulsc_mulb_ps46 & multm_reduce_mulsc_mulb_pc46;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy47 = multm_reduce_mulsc_mulb_ps47 & multm_reduce_mulsc_mulb_pc47;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy48 = multm_reduce_mulsc_mulb_ps48 & multm_reduce_mulsc_mulb_pc48;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy49 = multm_reduce_mulsc_mulb_ps49 & multm_reduce_mulsc_mulb_pc49;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy50 = multm_reduce_mulsc_mulb_ps50 & multm_reduce_mulsc_mulb_pc50;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy51 = multm_reduce_mulsc_mulb_ps51 & multm_reduce_mulsc_mulb_pc51;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy52 = multm_reduce_mulsc_mulb_ps52 & multm_reduce_mulsc_mulb_pc52;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy53 = multm_reduce_mulsc_mulb_ps53 & multm_reduce_mulsc_mulb_pc53;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy54 = multm_reduce_mulsc_mulb_ps54 & multm_reduce_mulsc_mulb_pc54;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy55 = multm_reduce_mulsc_mulb_ps55 & multm_reduce_mulsc_mulb_pc55;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy56 = multm_reduce_mulsc_mulb_ps56 & multm_reduce_mulsc_mulb_pc56;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy57 = multm_reduce_mulsc_mulb_ps57 & multm_reduce_mulsc_mulb_pc57;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy58 = multm_reduce_mulsc_mulb_ps58 & multm_reduce_mulsc_mulb_pc58;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy59 = multm_reduce_mulsc_mulb_ps59 & multm_reduce_mulsc_mulb_pc59;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy60 = multm_reduce_mulsc_mulb_ps60 & multm_reduce_mulsc_mulb_pc60;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy61 = multm_reduce_mulsc_mulb_ps61 & multm_reduce_mulsc_mulb_pc61;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy62 = multm_reduce_mulsc_mulb_ps62 & multm_reduce_mulsc_mulb_pc62;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy63 = multm_reduce_mulsc_mulb_ps63 & multm_reduce_mulsc_mulb_pc63;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy64 = multm_reduce_mulsc_mulb_ps64 & multm_reduce_mulsc_mulb_pc64;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy65 = multm_reduce_mulsc_mulb_ps65 & multm_reduce_mulsc_mulb_pc65;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy66 = multm_reduce_mulsc_mulb_ps66 & multm_reduce_mulsc_mulb_pc66;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy67 = multm_reduce_mulsc_mulb_ps67 & multm_reduce_mulsc_mulb_pc67;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy68 = multm_reduce_mulsc_mulb_ps68 & multm_reduce_mulsc_mulb_pc68;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy69 = multm_reduce_mulsc_mulb_ps69 & multm_reduce_mulsc_mulb_pc69;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy70 = multm_reduce_mulsc_mulb_ps70 & multm_reduce_mulsc_mulb_pc70;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy71 = multm_reduce_mulsc_mulb_ps71 & multm_reduce_mulsc_mulb_pc71;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy72 = multm_reduce_mulsc_mulb_ps72 & multm_reduce_mulsc_mulb_pc72;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy73 = multm_reduce_mulsc_mulb_ps73 & multm_reduce_mulsc_mulb_pc73;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy74 = multm_reduce_mulsc_mulb_ps74 & multm_reduce_mulsc_mulb_pc74;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy75 = multm_reduce_mulsc_mulb_ps75 & multm_reduce_mulsc_mulb_pc75;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy76 = multm_reduce_mulsc_mulb_ps76 & multm_reduce_mulsc_mulb_pc76;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy77 = multm_reduce_mulsc_mulb_ps77 & multm_reduce_mulsc_mulb_pc77;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy78 = multm_reduce_mulsc_mulb_ps78 & multm_reduce_mulsc_mulb_pc78;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy79 = multm_reduce_mulsc_mulb_ps79 & multm_reduce_mulsc_mulb_pc79;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy80 = multm_reduce_mulsc_mulb_ps80 & multm_reduce_mulsc_mulb_pc80;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy81 = multm_reduce_mulsc_mulb_ps81 & multm_reduce_mulsc_mulb_pc81;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy82 = multm_reduce_mulsc_mulb_ps82 & multm_reduce_mulsc_mulb_pc82;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy83 = multm_reduce_mulsc_mulb_ps83 & multm_reduce_mulsc_mulb_pc83;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy84 = multm_reduce_mulsc_mulb_ps84 & multm_reduce_mulsc_mulb_pc84;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy85 = multm_reduce_mulsc_mulb_ps85 & multm_reduce_mulsc_mulb_pc85;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy86 = multm_reduce_mulsc_mulb_ps86 & multm_reduce_mulsc_mulb_pc86;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy87 = multm_reduce_mulsc_mulb_ps87 & multm_reduce_mulsc_mulb_pc87;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy88 = multm_reduce_mulsc_mulb_ps88 & multm_reduce_mulsc_mulb_pc88;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy89 = multm_reduce_mulsc_mulb_ps89 & multm_reduce_mulsc_mulb_pc89;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy90 = multm_reduce_mulsc_mulb_ps90 & multm_reduce_mulsc_mulb_pc90;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy91 = multm_reduce_mulsc_mulb_ps91 & multm_reduce_mulsc_mulb_pc91;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy92 = multm_reduce_mulsc_mulb_ps92 & multm_reduce_mulsc_mulb_pc92;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy93 = multm_reduce_mulsc_mulb_ps93 & multm_reduce_mulsc_mulb_pc93;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy94 = multm_reduce_mulsc_mulb_ps94 & multm_reduce_mulsc_mulb_pc94;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy95 = multm_reduce_mulsc_mulb_ps95 & multm_reduce_mulsc_mulb_pc95;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy96 = multm_reduce_mulsc_mulb_ps96 & multm_reduce_mulsc_mulb_pc96;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy97 = multm_reduce_mulsc_mulb_ps97 & multm_reduce_mulsc_mulb_pc97;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy98 = multm_reduce_mulsc_mulb_ps98 & multm_reduce_mulsc_mulb_pc98;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy99 = multm_reduce_mulsc_mulb_ps99 & multm_reduce_mulsc_mulb_pc99;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy100 = multm_reduce_mulsc_mulb_ps100 & multm_reduce_mulsc_mulb_pc100;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy101 = multm_reduce_mulsc_mulb_ps101 & multm_reduce_mulsc_mulb_pc101;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy102 = multm_reduce_mulsc_mulb_ps102 & multm_reduce_mulsc_mulb_pc102;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy103 = multm_reduce_mulsc_mulb_ps103 & multm_reduce_mulsc_mulb_pc103;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy104 = multm_reduce_mulsc_mulb_ps104 & multm_reduce_mulsc_mulb_pc104;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy105 = multm_reduce_mulsc_mulb_ps105 & multm_reduce_mulsc_mulb_pc105;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy106 = multm_reduce_mulsc_mulb_ps106 & multm_reduce_mulsc_mulb_pc106;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy107 = multm_reduce_mulsc_mulb_ps107 & multm_reduce_mulsc_mulb_pc107;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy108 = multm_reduce_mulsc_mulb_ps108 & multm_reduce_mulsc_mulb_pc108;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy109 = multm_reduce_mulsc_mulb_ps109 & multm_reduce_mulsc_mulb_pc109;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy110 = multm_reduce_mulsc_mulb_ps110 & multm_reduce_mulsc_mulb_pc110;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy111 = multm_reduce_mulsc_mulb_ps111 & multm_reduce_mulsc_mulb_pc111;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy112 = multm_reduce_mulsc_mulb_ps112 & multm_reduce_mulsc_mulb_pc112;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy113 = multm_reduce_mulsc_mulb_ps113 & multm_reduce_mulsc_mulb_pc113;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy114 = multm_reduce_mulsc_mulb_ps114 & multm_reduce_mulsc_mulb_pc114;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy115 = multm_reduce_mulsc_mulb_ps115 & multm_reduce_mulsc_mulb_pc115;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy116 = multm_reduce_mulsc_mulb_ps116 & multm_reduce_mulsc_mulb_pc116;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy117 = multm_reduce_mulsc_mulb_ps117 & multm_reduce_mulsc_mulb_pc117;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy118 = multm_reduce_mulsc_mulb_ps118 & multm_reduce_mulsc_mulb_pc118;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy119 = multm_reduce_mulsc_mulb_ps119 & multm_reduce_mulsc_mulb_pc119;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy120 = multm_reduce_mulsc_mulb_ps120 & multm_reduce_mulsc_mulb_pc120;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy121 = multm_reduce_mulsc_mulb_ps121 & multm_reduce_mulsc_mulb_pc121;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy122 = multm_reduce_mulsc_mulb_ps122 & multm_reduce_mulsc_mulb_pc122;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy123 = multm_reduce_mulsc_mulb_ps123 & multm_reduce_mulsc_mulb_pc123;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy124 = multm_reduce_mulsc_mulb_ps124 & multm_reduce_mulsc_mulb_pc124;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy125 = multm_reduce_mulsc_mulb_ps125 & multm_reduce_mulsc_mulb_pc125;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy126 = multm_reduce_mulsc_mulb_ps126 & multm_reduce_mulsc_mulb_pc126;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy127 = multm_reduce_mulsc_mulb_ps127 & multm_reduce_mulsc_mulb_pc127;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy128 = multm_reduce_mulsc_mulb_ps128 & multm_reduce_mulsc_mulb_pc128;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy129 = multm_reduce_mulsc_mulb_ps129 & multm_reduce_mulsc_mulb_pc129;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy130 = multm_reduce_mulsc_mulb_ps130 & multm_reduce_mulsc_mulb_pc130;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy131 = multm_reduce_mulsc_mulb_ps131 & multm_reduce_mulsc_mulb_pc131;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy132 = multm_reduce_mulsc_mulb_ps132 & multm_reduce_mulsc_mulb_pc132;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy133 = multm_reduce_mulsc_mulb_ps133 & multm_reduce_mulsc_mulb_pc133;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy134 = multm_reduce_mulsc_mulb_ps134 & multm_reduce_mulsc_mulb_pc134;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy135 = multm_reduce_mulsc_mulb_ps135 & multm_reduce_mulsc_mulb_pc135;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy136 = multm_reduce_mulsc_mulb_ps136 & multm_reduce_mulsc_mulb_pc136;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy137 = multm_reduce_mulsc_mulb_ps137 & multm_reduce_mulsc_mulb_pc137;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy138 = multm_reduce_mulsc_mulb_ps138 & multm_reduce_mulsc_mulb_pc138;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy139 = multm_reduce_mulsc_mulb_ps139 & multm_reduce_mulsc_mulb_pc139;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy140 = multm_reduce_mulsc_mulb_ps140 & multm_reduce_mulsc_mulb_pc140;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy141 = multm_reduce_mulsc_mulb_ps141 & multm_reduce_mulsc_mulb_pc141;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy142 = multm_reduce_mulsc_mulb_ps142 & multm_reduce_mulsc_mulb_pc142;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy143 = multm_reduce_mulsc_mulb_ps143 & multm_reduce_mulsc_mulb_pc143;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy144 = multm_reduce_mulsc_mulb_ps144 & multm_reduce_mulsc_mulb_pc144;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy145 = multm_reduce_mulsc_mulb_ps145 & multm_reduce_mulsc_mulb_pc145;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy146 = multm_reduce_mulsc_mulb_ps146 & multm_reduce_mulsc_mulb_pc146;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy147 = multm_reduce_mulsc_mulb_ps147 & multm_reduce_mulsc_mulb_pc147;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy148 = multm_reduce_mulsc_mulb_ps148 & multm_reduce_mulsc_mulb_pc148;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy149 = multm_reduce_mulsc_mulb_ps149 & multm_reduce_mulsc_mulb_pc149;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy150 = multm_reduce_mulsc_mulb_ps150 & multm_reduce_mulsc_mulb_pc150;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy151 = multm_reduce_mulsc_mulb_ps151 & multm_reduce_mulsc_mulb_pc151;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy152 = multm_reduce_mulsc_mulb_ps152 & multm_reduce_mulsc_mulb_pc152;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy153 = multm_reduce_mulsc_mulb_ps153 & multm_reduce_mulsc_mulb_pc153;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy154 = multm_reduce_mulsc_mulb_ps154 & multm_reduce_mulsc_mulb_pc154;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy155 = multm_reduce_mulsc_mulb_ps155 & multm_reduce_mulsc_mulb_pc155;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy156 = multm_reduce_mulsc_mulb_ps156 & multm_reduce_mulsc_mulb_pc156;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy157 = multm_reduce_mulsc_mulb_ps157 & multm_reduce_mulsc_mulb_pc157;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy158 = multm_reduce_mulsc_mulb_ps158 & multm_reduce_mulsc_mulb_pc158;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy159 = multm_reduce_mulsc_mulb_ps159 & multm_reduce_mulsc_mulb_pc159;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy160 = multm_reduce_mulsc_mulb_ps160 & multm_reduce_mulsc_mulb_pc160;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy161 = multm_reduce_mulsc_mulb_ps161 & multm_reduce_mulsc_mulb_pc161;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy162 = multm_reduce_mulsc_mulb_ps162 & multm_reduce_mulsc_mulb_pc162;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy163 = multm_reduce_mulsc_mulb_ps163 & multm_reduce_mulsc_mulb_pc163;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy164 = multm_reduce_mulsc_mulb_ps164 & multm_reduce_mulsc_mulb_pc164;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy165 = multm_reduce_mulsc_mulb_ps165 & multm_reduce_mulsc_mulb_pc165;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy166 = multm_reduce_mulsc_mulb_ps166 & multm_reduce_mulsc_mulb_pc166;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy167 = multm_reduce_mulsc_mulb_ps167 & multm_reduce_mulsc_mulb_pc167;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy168 = multm_reduce_mulsc_mulb_ps168 & multm_reduce_mulsc_mulb_pc168;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy169 = multm_reduce_mulsc_mulb_ps169 & multm_reduce_mulsc_mulb_pc169;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy170 = multm_reduce_mulsc_mulb_ps170 & multm_reduce_mulsc_mulb_pc170;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy171 = multm_reduce_mulsc_mulb_ps171 & multm_reduce_mulsc_mulb_pc171;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy172 = multm_reduce_mulsc_mulb_ps172 & multm_reduce_mulsc_mulb_pc172;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy173 = multm_reduce_mulsc_mulb_ps173 & multm_reduce_mulsc_mulb_pc173;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy174 = multm_reduce_mulsc_mulb_ps174 & multm_reduce_mulsc_mulb_pc174;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy175 = multm_reduce_mulsc_mulb_ps175 & multm_reduce_mulsc_mulb_pc175;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy176 = multm_reduce_mulsc_mulb_ps176 & multm_reduce_mulsc_mulb_pc176;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy177 = multm_reduce_mulsc_mulb_ps177 & multm_reduce_mulsc_mulb_pc177;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy178 = multm_reduce_mulsc_mulb_ps178 & multm_reduce_mulsc_mulb_pc178;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy179 = multm_reduce_mulsc_mulb_ps179 & multm_reduce_mulsc_mulb_pc179;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy180 = multm_reduce_mulsc_mulb_ps180 & multm_reduce_mulsc_mulb_pc180;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy181 = multm_reduce_mulsc_mulb_ps181 & multm_reduce_mulsc_mulb_pc181;
  assign multm_reduce_mulsc_mulb_add3b1_maj3b_xy182 = multm_reduce_mulsc_mulb_ps182 & multm_reduce_mulsc_mulb_pc182;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx0 = multm_reduce_mulsc_mulb_yoc0 ^ multm_reduce_mulsc_mulb_ps0;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx1 = multm_reduce_mulsc_mulb_yoc1 ^ multm_reduce_mulsc_mulb_ps1;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx2 = multm_reduce_mulsc_mulb_yoc2 ^ multm_reduce_mulsc_mulb_ps2;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx3 = multm_reduce_mulsc_mulb_yoc3 ^ multm_reduce_mulsc_mulb_ps3;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx4 = multm_reduce_mulsc_mulb_yoc4 ^ multm_reduce_mulsc_mulb_ps4;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx5 = multm_reduce_mulsc_mulb_yoc5 ^ multm_reduce_mulsc_mulb_ps5;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx6 = multm_reduce_mulsc_mulb_yoc6 ^ multm_reduce_mulsc_mulb_ps6;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx7 = multm_reduce_mulsc_mulb_yoc7 ^ multm_reduce_mulsc_mulb_ps7;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx8 = multm_reduce_mulsc_mulb_yoc8 ^ multm_reduce_mulsc_mulb_ps8;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx9 = multm_reduce_mulsc_mulb_yoc9 ^ multm_reduce_mulsc_mulb_ps9;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx10 = multm_reduce_mulsc_mulb_yoc10 ^ multm_reduce_mulsc_mulb_ps10;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx11 = multm_reduce_mulsc_mulb_yoc11 ^ multm_reduce_mulsc_mulb_ps11;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx12 = multm_reduce_mulsc_mulb_yoc12 ^ multm_reduce_mulsc_mulb_ps12;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx13 = multm_reduce_mulsc_mulb_yoc13 ^ multm_reduce_mulsc_mulb_ps13;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx14 = multm_reduce_mulsc_mulb_yoc14 ^ multm_reduce_mulsc_mulb_ps14;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx15 = multm_reduce_mulsc_mulb_yoc15 ^ multm_reduce_mulsc_mulb_ps15;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx16 = multm_reduce_mulsc_mulb_yoc16 ^ multm_reduce_mulsc_mulb_ps16;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx17 = multm_reduce_mulsc_mulb_yoc17 ^ multm_reduce_mulsc_mulb_ps17;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx18 = multm_reduce_mulsc_mulb_yoc18 ^ multm_reduce_mulsc_mulb_ps18;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx19 = multm_reduce_mulsc_mulb_yoc19 ^ multm_reduce_mulsc_mulb_ps19;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx20 = multm_reduce_mulsc_mulb_yoc20 ^ multm_reduce_mulsc_mulb_ps20;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx21 = multm_reduce_mulsc_mulb_yoc21 ^ multm_reduce_mulsc_mulb_ps21;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx22 = multm_reduce_mulsc_mulb_yoc22 ^ multm_reduce_mulsc_mulb_ps22;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx23 = multm_reduce_mulsc_mulb_yoc23 ^ multm_reduce_mulsc_mulb_ps23;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx24 = multm_reduce_mulsc_mulb_yoc24 ^ multm_reduce_mulsc_mulb_ps24;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx25 = multm_reduce_mulsc_mulb_yoc25 ^ multm_reduce_mulsc_mulb_ps25;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx26 = multm_reduce_mulsc_mulb_yoc26 ^ multm_reduce_mulsc_mulb_ps26;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx27 = multm_reduce_mulsc_mulb_yoc27 ^ multm_reduce_mulsc_mulb_ps27;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx28 = multm_reduce_mulsc_mulb_yoc28 ^ multm_reduce_mulsc_mulb_ps28;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx29 = multm_reduce_mulsc_mulb_yoc29 ^ multm_reduce_mulsc_mulb_ps29;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx30 = multm_reduce_mulsc_mulb_yoc30 ^ multm_reduce_mulsc_mulb_ps30;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx31 = multm_reduce_mulsc_mulb_yoc31 ^ multm_reduce_mulsc_mulb_ps31;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx32 = multm_reduce_mulsc_mulb_yoc32 ^ multm_reduce_mulsc_mulb_ps32;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx33 = multm_reduce_mulsc_mulb_yoc33 ^ multm_reduce_mulsc_mulb_ps33;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx34 = multm_reduce_mulsc_mulb_yoc34 ^ multm_reduce_mulsc_mulb_ps34;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx35 = multm_reduce_mulsc_mulb_yoc35 ^ multm_reduce_mulsc_mulb_ps35;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx36 = multm_reduce_mulsc_mulb_yoc36 ^ multm_reduce_mulsc_mulb_ps36;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx37 = multm_reduce_mulsc_mulb_yoc37 ^ multm_reduce_mulsc_mulb_ps37;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx38 = multm_reduce_mulsc_mulb_yoc38 ^ multm_reduce_mulsc_mulb_ps38;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx39 = multm_reduce_mulsc_mulb_yoc39 ^ multm_reduce_mulsc_mulb_ps39;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx40 = multm_reduce_mulsc_mulb_yoc40 ^ multm_reduce_mulsc_mulb_ps40;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx41 = multm_reduce_mulsc_mulb_yoc41 ^ multm_reduce_mulsc_mulb_ps41;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx42 = multm_reduce_mulsc_mulb_yoc42 ^ multm_reduce_mulsc_mulb_ps42;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx43 = multm_reduce_mulsc_mulb_yoc43 ^ multm_reduce_mulsc_mulb_ps43;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx44 = multm_reduce_mulsc_mulb_yoc44 ^ multm_reduce_mulsc_mulb_ps44;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx45 = multm_reduce_mulsc_mulb_yoc45 ^ multm_reduce_mulsc_mulb_ps45;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx46 = multm_reduce_mulsc_mulb_yoc46 ^ multm_reduce_mulsc_mulb_ps46;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx47 = multm_reduce_mulsc_mulb_yoc47 ^ multm_reduce_mulsc_mulb_ps47;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx48 = multm_reduce_mulsc_mulb_yoc48 ^ multm_reduce_mulsc_mulb_ps48;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx49 = multm_reduce_mulsc_mulb_yoc49 ^ multm_reduce_mulsc_mulb_ps49;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx50 = multm_reduce_mulsc_mulb_yoc50 ^ multm_reduce_mulsc_mulb_ps50;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx51 = multm_reduce_mulsc_mulb_yoc51 ^ multm_reduce_mulsc_mulb_ps51;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx52 = multm_reduce_mulsc_mulb_yoc52 ^ multm_reduce_mulsc_mulb_ps52;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx53 = multm_reduce_mulsc_mulb_yoc53 ^ multm_reduce_mulsc_mulb_ps53;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx54 = multm_reduce_mulsc_mulb_yoc54 ^ multm_reduce_mulsc_mulb_ps54;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx55 = multm_reduce_mulsc_mulb_yoc55 ^ multm_reduce_mulsc_mulb_ps55;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx56 = multm_reduce_mulsc_mulb_yoc56 ^ multm_reduce_mulsc_mulb_ps56;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx57 = multm_reduce_mulsc_mulb_yoc57 ^ multm_reduce_mulsc_mulb_ps57;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx58 = multm_reduce_mulsc_mulb_yoc58 ^ multm_reduce_mulsc_mulb_ps58;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx59 = multm_reduce_mulsc_mulb_yoc59 ^ multm_reduce_mulsc_mulb_ps59;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx60 = multm_reduce_mulsc_mulb_yoc60 ^ multm_reduce_mulsc_mulb_ps60;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx61 = multm_reduce_mulsc_mulb_yoc61 ^ multm_reduce_mulsc_mulb_ps61;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx62 = multm_reduce_mulsc_mulb_yoc62 ^ multm_reduce_mulsc_mulb_ps62;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx63 = multm_reduce_mulsc_mulb_yoc63 ^ multm_reduce_mulsc_mulb_ps63;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx64 = multm_reduce_mulsc_mulb_yoc64 ^ multm_reduce_mulsc_mulb_ps64;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx65 = multm_reduce_mulsc_mulb_yoc65 ^ multm_reduce_mulsc_mulb_ps65;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx66 = multm_reduce_mulsc_mulb_yoc66 ^ multm_reduce_mulsc_mulb_ps66;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx67 = multm_reduce_mulsc_mulb_yoc67 ^ multm_reduce_mulsc_mulb_ps67;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx68 = multm_reduce_mulsc_mulb_yoc68 ^ multm_reduce_mulsc_mulb_ps68;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx69 = multm_reduce_mulsc_mulb_yoc69 ^ multm_reduce_mulsc_mulb_ps69;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx70 = multm_reduce_mulsc_mulb_yoc70 ^ multm_reduce_mulsc_mulb_ps70;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx71 = multm_reduce_mulsc_mulb_yoc71 ^ multm_reduce_mulsc_mulb_ps71;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx72 = multm_reduce_mulsc_mulb_yoc72 ^ multm_reduce_mulsc_mulb_ps72;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx73 = multm_reduce_mulsc_mulb_yoc73 ^ multm_reduce_mulsc_mulb_ps73;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx74 = multm_reduce_mulsc_mulb_yoc74 ^ multm_reduce_mulsc_mulb_ps74;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx75 = multm_reduce_mulsc_mulb_yoc75 ^ multm_reduce_mulsc_mulb_ps75;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx76 = multm_reduce_mulsc_mulb_yoc76 ^ multm_reduce_mulsc_mulb_ps76;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx77 = multm_reduce_mulsc_mulb_yoc77 ^ multm_reduce_mulsc_mulb_ps77;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx78 = multm_reduce_mulsc_mulb_yoc78 ^ multm_reduce_mulsc_mulb_ps78;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx79 = multm_reduce_mulsc_mulb_yoc79 ^ multm_reduce_mulsc_mulb_ps79;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx80 = multm_reduce_mulsc_mulb_yoc80 ^ multm_reduce_mulsc_mulb_ps80;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx81 = multm_reduce_mulsc_mulb_yoc81 ^ multm_reduce_mulsc_mulb_ps81;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx82 = multm_reduce_mulsc_mulb_yoc82 ^ multm_reduce_mulsc_mulb_ps82;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx83 = multm_reduce_mulsc_mulb_yoc83 ^ multm_reduce_mulsc_mulb_ps83;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx84 = multm_reduce_mulsc_mulb_yoc84 ^ multm_reduce_mulsc_mulb_ps84;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx85 = multm_reduce_mulsc_mulb_yoc85 ^ multm_reduce_mulsc_mulb_ps85;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx86 = multm_reduce_mulsc_mulb_yoc86 ^ multm_reduce_mulsc_mulb_ps86;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx87 = multm_reduce_mulsc_mulb_yoc87 ^ multm_reduce_mulsc_mulb_ps87;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx88 = multm_reduce_mulsc_mulb_yoc88 ^ multm_reduce_mulsc_mulb_ps88;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx89 = multm_reduce_mulsc_mulb_yoc89 ^ multm_reduce_mulsc_mulb_ps89;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx90 = multm_reduce_mulsc_mulb_yoc90 ^ multm_reduce_mulsc_mulb_ps90;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx91 = multm_reduce_mulsc_mulb_yoc91 ^ multm_reduce_mulsc_mulb_ps91;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx92 = multm_reduce_mulsc_mulb_yoc92 ^ multm_reduce_mulsc_mulb_ps92;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx93 = multm_reduce_mulsc_mulb_yoc93 ^ multm_reduce_mulsc_mulb_ps93;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx94 = multm_reduce_mulsc_mulb_yoc94 ^ multm_reduce_mulsc_mulb_ps94;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx95 = multm_reduce_mulsc_mulb_yoc95 ^ multm_reduce_mulsc_mulb_ps95;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx96 = multm_reduce_mulsc_mulb_yoc96 ^ multm_reduce_mulsc_mulb_ps96;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx97 = multm_reduce_mulsc_mulb_yoc97 ^ multm_reduce_mulsc_mulb_ps97;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx98 = multm_reduce_mulsc_mulb_yoc98 ^ multm_reduce_mulsc_mulb_ps98;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx99 = multm_reduce_mulsc_mulb_yoc99 ^ multm_reduce_mulsc_mulb_ps99;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx100 = multm_reduce_mulsc_mulb_yoc100 ^ multm_reduce_mulsc_mulb_ps100;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx101 = multm_reduce_mulsc_mulb_yoc101 ^ multm_reduce_mulsc_mulb_ps101;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx102 = multm_reduce_mulsc_mulb_yoc102 ^ multm_reduce_mulsc_mulb_ps102;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx103 = multm_reduce_mulsc_mulb_yoc103 ^ multm_reduce_mulsc_mulb_ps103;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx104 = multm_reduce_mulsc_mulb_yoc104 ^ multm_reduce_mulsc_mulb_ps104;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx105 = multm_reduce_mulsc_mulb_yoc105 ^ multm_reduce_mulsc_mulb_ps105;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx106 = multm_reduce_mulsc_mulb_yoc106 ^ multm_reduce_mulsc_mulb_ps106;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx107 = multm_reduce_mulsc_mulb_yoc107 ^ multm_reduce_mulsc_mulb_ps107;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx108 = multm_reduce_mulsc_mulb_yoc108 ^ multm_reduce_mulsc_mulb_ps108;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx109 = multm_reduce_mulsc_mulb_yoc109 ^ multm_reduce_mulsc_mulb_ps109;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx110 = multm_reduce_mulsc_mulb_yoc110 ^ multm_reduce_mulsc_mulb_ps110;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx111 = multm_reduce_mulsc_mulb_yoc111 ^ multm_reduce_mulsc_mulb_ps111;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx112 = multm_reduce_mulsc_mulb_yoc112 ^ multm_reduce_mulsc_mulb_ps112;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx113 = multm_reduce_mulsc_mulb_yoc113 ^ multm_reduce_mulsc_mulb_ps113;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx114 = multm_reduce_mulsc_mulb_yoc114 ^ multm_reduce_mulsc_mulb_ps114;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx115 = multm_reduce_mulsc_mulb_yoc115 ^ multm_reduce_mulsc_mulb_ps115;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx116 = multm_reduce_mulsc_mulb_yoc116 ^ multm_reduce_mulsc_mulb_ps116;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx117 = multm_reduce_mulsc_mulb_yoc117 ^ multm_reduce_mulsc_mulb_ps117;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx118 = multm_reduce_mulsc_mulb_yoc118 ^ multm_reduce_mulsc_mulb_ps118;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx119 = multm_reduce_mulsc_mulb_yoc119 ^ multm_reduce_mulsc_mulb_ps119;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx120 = multm_reduce_mulsc_mulb_yoc120 ^ multm_reduce_mulsc_mulb_ps120;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx121 = multm_reduce_mulsc_mulb_yoc121 ^ multm_reduce_mulsc_mulb_ps121;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx122 = multm_reduce_mulsc_mulb_yoc122 ^ multm_reduce_mulsc_mulb_ps122;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx123 = multm_reduce_mulsc_mulb_yoc123 ^ multm_reduce_mulsc_mulb_ps123;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx124 = multm_reduce_mulsc_mulb_yoc124 ^ multm_reduce_mulsc_mulb_ps124;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx125 = multm_reduce_mulsc_mulb_yoc125 ^ multm_reduce_mulsc_mulb_ps125;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx126 = multm_reduce_mulsc_mulb_yoc126 ^ multm_reduce_mulsc_mulb_ps126;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx127 = multm_reduce_mulsc_mulb_yoc127 ^ multm_reduce_mulsc_mulb_ps127;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx128 = multm_reduce_mulsc_mulb_yoc128 ^ multm_reduce_mulsc_mulb_ps128;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx129 = multm_reduce_mulsc_mulb_yoc129 ^ multm_reduce_mulsc_mulb_ps129;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx130 = multm_reduce_mulsc_mulb_yoc130 ^ multm_reduce_mulsc_mulb_ps130;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx131 = multm_reduce_mulsc_mulb_yoc131 ^ multm_reduce_mulsc_mulb_ps131;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx132 = multm_reduce_mulsc_mulb_yoc132 ^ multm_reduce_mulsc_mulb_ps132;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx133 = multm_reduce_mulsc_mulb_yoc133 ^ multm_reduce_mulsc_mulb_ps133;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx134 = multm_reduce_mulsc_mulb_yoc134 ^ multm_reduce_mulsc_mulb_ps134;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx135 = multm_reduce_mulsc_mulb_yoc135 ^ multm_reduce_mulsc_mulb_ps135;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx136 = multm_reduce_mulsc_mulb_yoc136 ^ multm_reduce_mulsc_mulb_ps136;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx137 = multm_reduce_mulsc_mulb_yoc137 ^ multm_reduce_mulsc_mulb_ps137;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx138 = multm_reduce_mulsc_mulb_yoc138 ^ multm_reduce_mulsc_mulb_ps138;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx139 = multm_reduce_mulsc_mulb_yoc139 ^ multm_reduce_mulsc_mulb_ps139;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx140 = multm_reduce_mulsc_mulb_yoc140 ^ multm_reduce_mulsc_mulb_ps140;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx141 = multm_reduce_mulsc_mulb_yoc141 ^ multm_reduce_mulsc_mulb_ps141;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx142 = multm_reduce_mulsc_mulb_yoc142 ^ multm_reduce_mulsc_mulb_ps142;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx143 = multm_reduce_mulsc_mulb_yoc143 ^ multm_reduce_mulsc_mulb_ps143;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx144 = multm_reduce_mulsc_mulb_yoc144 ^ multm_reduce_mulsc_mulb_ps144;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx145 = multm_reduce_mulsc_mulb_yoc145 ^ multm_reduce_mulsc_mulb_ps145;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx146 = multm_reduce_mulsc_mulb_yoc146 ^ multm_reduce_mulsc_mulb_ps146;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx147 = multm_reduce_mulsc_mulb_yoc147 ^ multm_reduce_mulsc_mulb_ps147;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx148 = multm_reduce_mulsc_mulb_yoc148 ^ multm_reduce_mulsc_mulb_ps148;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx149 = multm_reduce_mulsc_mulb_yoc149 ^ multm_reduce_mulsc_mulb_ps149;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx150 = multm_reduce_mulsc_mulb_yoc150 ^ multm_reduce_mulsc_mulb_ps150;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx151 = multm_reduce_mulsc_mulb_yoc151 ^ multm_reduce_mulsc_mulb_ps151;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx152 = multm_reduce_mulsc_mulb_yoc152 ^ multm_reduce_mulsc_mulb_ps152;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx153 = multm_reduce_mulsc_mulb_yoc153 ^ multm_reduce_mulsc_mulb_ps153;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx154 = multm_reduce_mulsc_mulb_yoc154 ^ multm_reduce_mulsc_mulb_ps154;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx155 = multm_reduce_mulsc_mulb_yoc155 ^ multm_reduce_mulsc_mulb_ps155;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx156 = multm_reduce_mulsc_mulb_yoc156 ^ multm_reduce_mulsc_mulb_ps156;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx157 = multm_reduce_mulsc_mulb_yoc157 ^ multm_reduce_mulsc_mulb_ps157;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx158 = multm_reduce_mulsc_mulb_yoc158 ^ multm_reduce_mulsc_mulb_ps158;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx159 = multm_reduce_mulsc_mulb_yoc159 ^ multm_reduce_mulsc_mulb_ps159;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx160 = multm_reduce_mulsc_mulb_yoc160 ^ multm_reduce_mulsc_mulb_ps160;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx161 = multm_reduce_mulsc_mulb_yoc161 ^ multm_reduce_mulsc_mulb_ps161;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx162 = multm_reduce_mulsc_mulb_yoc162 ^ multm_reduce_mulsc_mulb_ps162;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx163 = multm_reduce_mulsc_mulb_yoc163 ^ multm_reduce_mulsc_mulb_ps163;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx164 = multm_reduce_mulsc_mulb_yoc164 ^ multm_reduce_mulsc_mulb_ps164;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx165 = multm_reduce_mulsc_mulb_yoc165 ^ multm_reduce_mulsc_mulb_ps165;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx166 = multm_reduce_mulsc_mulb_yoc166 ^ multm_reduce_mulsc_mulb_ps166;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx167 = multm_reduce_mulsc_mulb_yoc167 ^ multm_reduce_mulsc_mulb_ps167;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx168 = multm_reduce_mulsc_mulb_yoc168 ^ multm_reduce_mulsc_mulb_ps168;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx169 = multm_reduce_mulsc_mulb_yoc169 ^ multm_reduce_mulsc_mulb_ps169;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx170 = multm_reduce_mulsc_mulb_yoc170 ^ multm_reduce_mulsc_mulb_ps170;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx171 = multm_reduce_mulsc_mulb_yoc171 ^ multm_reduce_mulsc_mulb_ps171;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx172 = multm_reduce_mulsc_mulb_yoc172 ^ multm_reduce_mulsc_mulb_ps172;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx173 = multm_reduce_mulsc_mulb_yoc173 ^ multm_reduce_mulsc_mulb_ps173;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx174 = multm_reduce_mulsc_mulb_yoc174 ^ multm_reduce_mulsc_mulb_ps174;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx175 = multm_reduce_mulsc_mulb_yoc175 ^ multm_reduce_mulsc_mulb_ps175;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx176 = multm_reduce_mulsc_mulb_yoc176 ^ multm_reduce_mulsc_mulb_ps176;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx177 = multm_reduce_mulsc_mulb_yoc177 ^ multm_reduce_mulsc_mulb_ps177;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx178 = multm_reduce_mulsc_mulb_yoc178 ^ multm_reduce_mulsc_mulb_ps178;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx179 = multm_reduce_mulsc_mulb_yoc179 ^ multm_reduce_mulsc_mulb_ps179;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx180 = multm_reduce_mulsc_mulb_yoc180 ^ multm_reduce_mulsc_mulb_ps180;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx181 = multm_reduce_mulsc_mulb_yoc181 ^ multm_reduce_mulsc_mulb_ps181;
  assign multm_reduce_mulsc_mulb_add3b1_xor3b_wx182 = multm_reduce_mulsc_mulb_yoc182 ^ multm_reduce_mulsc_mulb_ps182;
  assign multm_reduce_mulsc_mulb_cq0 = xn3 & multm_reduce_sb0;
  assign multm_reduce_mulsc_mulb_cq1 = xn3 & multm_reduce_sb1;
  assign multm_reduce_mulsc_mulb_cq2 = xn3 & multm_reduce_sb2;
  assign multm_reduce_mulsc_mulb_cq3 = xn3 & multm_reduce_sb3;
  assign multm_reduce_mulsc_mulb_cq4 = xn3 & multm_reduce_sb4;
  assign multm_reduce_mulsc_mulb_cq5 = xn3 & multm_reduce_sb5;
  assign multm_reduce_mulsc_mulb_cq6 = xn3 & multm_reduce_sb6;
  assign multm_reduce_mulsc_mulb_cq7 = xn3 & multm_reduce_sb7;
  assign multm_reduce_mulsc_mulb_cq8 = xn3 & multm_reduce_sb8;
  assign multm_reduce_mulsc_mulb_cq9 = xn3 & multm_reduce_sb9;
  assign multm_reduce_mulsc_mulb_cq10 = xn3 & multm_reduce_sb10;
  assign multm_reduce_mulsc_mulb_cq11 = xn3 & multm_reduce_sb11;
  assign multm_reduce_mulsc_mulb_cq12 = xn3 & multm_reduce_sb12;
  assign multm_reduce_mulsc_mulb_cq13 = xn3 & multm_reduce_sb13;
  assign multm_reduce_mulsc_mulb_cq14 = xn3 & multm_reduce_sb14;
  assign multm_reduce_mulsc_mulb_cq15 = xn3 & multm_reduce_sb15;
  assign multm_reduce_mulsc_mulb_cq16 = xn3 & multm_reduce_sb16;
  assign multm_reduce_mulsc_mulb_cq17 = xn3 & multm_reduce_sb17;
  assign multm_reduce_mulsc_mulb_cq18 = xn3 & multm_reduce_sb18;
  assign multm_reduce_mulsc_mulb_cq19 = xn3 & multm_reduce_sb19;
  assign multm_reduce_mulsc_mulb_cq20 = xn3 & multm_reduce_sb20;
  assign multm_reduce_mulsc_mulb_cq21 = xn3 & multm_reduce_sb21;
  assign multm_reduce_mulsc_mulb_cq22 = xn3 & multm_reduce_sb22;
  assign multm_reduce_mulsc_mulb_cq23 = xn3 & multm_reduce_sb23;
  assign multm_reduce_mulsc_mulb_cq24 = xn3 & multm_reduce_sb24;
  assign multm_reduce_mulsc_mulb_cq25 = xn3 & multm_reduce_sb25;
  assign multm_reduce_mulsc_mulb_cq26 = xn3 & multm_reduce_sb26;
  assign multm_reduce_mulsc_mulb_cq27 = xn3 & multm_reduce_sb27;
  assign multm_reduce_mulsc_mulb_cq28 = xn3 & multm_reduce_sb28;
  assign multm_reduce_mulsc_mulb_cq29 = xn3 & multm_reduce_sb29;
  assign multm_reduce_mulsc_mulb_cq30 = xn3 & multm_reduce_sb30;
  assign multm_reduce_mulsc_mulb_cq31 = xn3 & multm_reduce_sb31;
  assign multm_reduce_mulsc_mulb_cq32 = xn3 & multm_reduce_sb32;
  assign multm_reduce_mulsc_mulb_cq33 = xn3 & multm_reduce_sb33;
  assign multm_reduce_mulsc_mulb_cq34 = xn3 & multm_reduce_sb34;
  assign multm_reduce_mulsc_mulb_cq35 = xn3 & multm_reduce_sb35;
  assign multm_reduce_mulsc_mulb_cq36 = xn3 & multm_reduce_sb36;
  assign multm_reduce_mulsc_mulb_cq37 = xn3 & multm_reduce_sb37;
  assign multm_reduce_mulsc_mulb_cq38 = xn3 & multm_reduce_sb38;
  assign multm_reduce_mulsc_mulb_cq39 = xn3 & multm_reduce_sb39;
  assign multm_reduce_mulsc_mulb_cq40 = xn3 & multm_reduce_sb40;
  assign multm_reduce_mulsc_mulb_cq41 = xn3 & multm_reduce_sb41;
  assign multm_reduce_mulsc_mulb_cq42 = xn3 & multm_reduce_sb42;
  assign multm_reduce_mulsc_mulb_cq43 = xn3 & multm_reduce_sb43;
  assign multm_reduce_mulsc_mulb_cq44 = xn3 & multm_reduce_sb44;
  assign multm_reduce_mulsc_mulb_cq45 = xn3 & multm_reduce_sb45;
  assign multm_reduce_mulsc_mulb_cq46 = xn3 & multm_reduce_sb46;
  assign multm_reduce_mulsc_mulb_cq47 = xn3 & multm_reduce_sb47;
  assign multm_reduce_mulsc_mulb_cq48 = xn3 & multm_reduce_sb48;
  assign multm_reduce_mulsc_mulb_cq49 = xn3 & multm_reduce_sb49;
  assign multm_reduce_mulsc_mulb_cq50 = xn3 & multm_reduce_sb50;
  assign multm_reduce_mulsc_mulb_cq51 = xn3 & multm_reduce_sb51;
  assign multm_reduce_mulsc_mulb_cq52 = xn3 & multm_reduce_sb52;
  assign multm_reduce_mulsc_mulb_cq53 = xn3 & multm_reduce_sb53;
  assign multm_reduce_mulsc_mulb_cq54 = xn3 & multm_reduce_sb54;
  assign multm_reduce_mulsc_mulb_cq55 = xn3 & multm_reduce_sb55;
  assign multm_reduce_mulsc_mulb_cq56 = xn3 & multm_reduce_sb56;
  assign multm_reduce_mulsc_mulb_cq57 = xn3 & multm_reduce_sb57;
  assign multm_reduce_mulsc_mulb_cq58 = xn3 & multm_reduce_sb58;
  assign multm_reduce_mulsc_mulb_cq59 = xn3 & multm_reduce_sb59;
  assign multm_reduce_mulsc_mulb_cq60 = xn3 & multm_reduce_sb60;
  assign multm_reduce_mulsc_mulb_cq61 = xn3 & multm_reduce_sb61;
  assign multm_reduce_mulsc_mulb_cq62 = xn3 & multm_reduce_sb62;
  assign multm_reduce_mulsc_mulb_cq63 = xn3 & multm_reduce_sb63;
  assign multm_reduce_mulsc_mulb_cq64 = xn3 & multm_reduce_sb64;
  assign multm_reduce_mulsc_mulb_cq65 = xn3 & multm_reduce_sb65;
  assign multm_reduce_mulsc_mulb_cq66 = xn3 & multm_reduce_sb66;
  assign multm_reduce_mulsc_mulb_cq67 = xn3 & multm_reduce_sb67;
  assign multm_reduce_mulsc_mulb_cq68 = xn3 & multm_reduce_sb68;
  assign multm_reduce_mulsc_mulb_cq69 = xn3 & multm_reduce_sb69;
  assign multm_reduce_mulsc_mulb_cq70 = xn3 & multm_reduce_sb70;
  assign multm_reduce_mulsc_mulb_cq71 = xn3 & multm_reduce_sb71;
  assign multm_reduce_mulsc_mulb_cq72 = xn3 & multm_reduce_sb72;
  assign multm_reduce_mulsc_mulb_cq73 = xn3 & multm_reduce_sb73;
  assign multm_reduce_mulsc_mulb_cq74 = xn3 & multm_reduce_sb74;
  assign multm_reduce_mulsc_mulb_cq75 = xn3 & multm_reduce_sb75;
  assign multm_reduce_mulsc_mulb_cq76 = xn3 & multm_reduce_sb76;
  assign multm_reduce_mulsc_mulb_cq77 = xn3 & multm_reduce_sb77;
  assign multm_reduce_mulsc_mulb_cq78 = xn3 & multm_reduce_sb78;
  assign multm_reduce_mulsc_mulb_cq79 = xn3 & multm_reduce_sb79;
  assign multm_reduce_mulsc_mulb_cq80 = xn3 & multm_reduce_sb80;
  assign multm_reduce_mulsc_mulb_cq81 = xn3 & multm_reduce_sb81;
  assign multm_reduce_mulsc_mulb_cq82 = xn3 & multm_reduce_sb82;
  assign multm_reduce_mulsc_mulb_cq83 = xn3 & multm_reduce_sb83;
  assign multm_reduce_mulsc_mulb_cq84 = xn3 & multm_reduce_sb84;
  assign multm_reduce_mulsc_mulb_cq85 = xn3 & multm_reduce_sb85;
  assign multm_reduce_mulsc_mulb_cq86 = xn3 & multm_reduce_sb86;
  assign multm_reduce_mulsc_mulb_cq87 = xn3 & multm_reduce_sb87;
  assign multm_reduce_mulsc_mulb_cq88 = xn3 & multm_reduce_sb88;
  assign multm_reduce_mulsc_mulb_cq89 = xn3 & multm_reduce_sb89;
  assign multm_reduce_mulsc_mulb_cq90 = xn3 & multm_reduce_sb90;
  assign multm_reduce_mulsc_mulb_cq91 = xn3 & multm_reduce_sb91;
  assign multm_reduce_mulsc_mulb_cq92 = xn3 & multm_reduce_sb92;
  assign multm_reduce_mulsc_mulb_cq93 = xn3 & multm_reduce_sb93;
  assign multm_reduce_mulsc_mulb_cq94 = xn3 & multm_reduce_sb94;
  assign multm_reduce_mulsc_mulb_cq95 = xn3 & multm_reduce_sb95;
  assign multm_reduce_mulsc_mulb_cq96 = xn3 & multm_reduce_sb96;
  assign multm_reduce_mulsc_mulb_cq97 = xn3 & multm_reduce_sb97;
  assign multm_reduce_mulsc_mulb_cq98 = xn3 & multm_reduce_sb98;
  assign multm_reduce_mulsc_mulb_cq99 = xn3 & multm_reduce_sb99;
  assign multm_reduce_mulsc_mulb_cq100 = xn3 & multm_reduce_sb100;
  assign multm_reduce_mulsc_mulb_cq101 = xn3 & multm_reduce_sb101;
  assign multm_reduce_mulsc_mulb_cq102 = xn3 & multm_reduce_sb102;
  assign multm_reduce_mulsc_mulb_cq103 = xn3 & multm_reduce_sb103;
  assign multm_reduce_mulsc_mulb_cq104 = xn3 & multm_reduce_sb104;
  assign multm_reduce_mulsc_mulb_cq105 = xn3 & multm_reduce_sb105;
  assign multm_reduce_mulsc_mulb_cq106 = xn3 & multm_reduce_sb106;
  assign multm_reduce_mulsc_mulb_cq107 = xn3 & multm_reduce_sb107;
  assign multm_reduce_mulsc_mulb_cq108 = xn3 & multm_reduce_sb108;
  assign multm_reduce_mulsc_mulb_cq109 = xn3 & multm_reduce_sb109;
  assign multm_reduce_mulsc_mulb_cq110 = xn3 & multm_reduce_sb110;
  assign multm_reduce_mulsc_mulb_cq111 = xn3 & multm_reduce_sb111;
  assign multm_reduce_mulsc_mulb_cq112 = xn3 & multm_reduce_sb112;
  assign multm_reduce_mulsc_mulb_cq113 = xn3 & multm_reduce_sb113;
  assign multm_reduce_mulsc_mulb_cq114 = xn3 & multm_reduce_sb114;
  assign multm_reduce_mulsc_mulb_cq115 = xn3 & multm_reduce_sb115;
  assign multm_reduce_mulsc_mulb_cq116 = xn3 & multm_reduce_sb116;
  assign multm_reduce_mulsc_mulb_cq117 = xn3 & multm_reduce_sb117;
  assign multm_reduce_mulsc_mulb_cq118 = xn3 & multm_reduce_sb118;
  assign multm_reduce_mulsc_mulb_cq119 = xn3 & multm_reduce_sb119;
  assign multm_reduce_mulsc_mulb_cq120 = xn3 & multm_reduce_sb120;
  assign multm_reduce_mulsc_mulb_cq121 = xn3 & multm_reduce_sb121;
  assign multm_reduce_mulsc_mulb_cq122 = xn3 & multm_reduce_sb122;
  assign multm_reduce_mulsc_mulb_cq123 = xn3 & multm_reduce_sb123;
  assign multm_reduce_mulsc_mulb_cq124 = xn3 & multm_reduce_sb124;
  assign multm_reduce_mulsc_mulb_cq125 = xn3 & multm_reduce_sb125;
  assign multm_reduce_mulsc_mulb_cq126 = xn3 & multm_reduce_sb126;
  assign multm_reduce_mulsc_mulb_cq127 = xn3 & multm_reduce_sb127;
  assign multm_reduce_mulsc_mulb_cq128 = xn3 & multm_reduce_sb128;
  assign multm_reduce_mulsc_mulb_cq129 = xn3 & multm_reduce_sb129;
  assign multm_reduce_mulsc_mulb_cq130 = xn3 & multm_reduce_sb130;
  assign multm_reduce_mulsc_mulb_cq131 = xn3 & multm_reduce_sb131;
  assign multm_reduce_mulsc_mulb_cq132 = xn3 & multm_reduce_sb132;
  assign multm_reduce_mulsc_mulb_cq133 = xn3 & multm_reduce_sb133;
  assign multm_reduce_mulsc_mulb_cq134 = xn3 & multm_reduce_sb134;
  assign multm_reduce_mulsc_mulb_cq135 = xn3 & multm_reduce_sb135;
  assign multm_reduce_mulsc_mulb_cq136 = xn3 & multm_reduce_sb136;
  assign multm_reduce_mulsc_mulb_cq137 = xn3 & multm_reduce_sb137;
  assign multm_reduce_mulsc_mulb_cq138 = xn3 & multm_reduce_sb138;
  assign multm_reduce_mulsc_mulb_cq139 = xn3 & multm_reduce_sb139;
  assign multm_reduce_mulsc_mulb_cq140 = xn3 & multm_reduce_sb140;
  assign multm_reduce_mulsc_mulb_cq141 = xn3 & multm_reduce_sb141;
  assign multm_reduce_mulsc_mulb_cq142 = xn3 & multm_reduce_sb142;
  assign multm_reduce_mulsc_mulb_cq143 = xn3 & multm_reduce_sb143;
  assign multm_reduce_mulsc_mulb_cq144 = xn3 & multm_reduce_sb144;
  assign multm_reduce_mulsc_mulb_cq145 = xn3 & multm_reduce_sb145;
  assign multm_reduce_mulsc_mulb_cq146 = xn3 & multm_reduce_sb146;
  assign multm_reduce_mulsc_mulb_cq147 = xn3 & multm_reduce_sb147;
  assign multm_reduce_mulsc_mulb_cq148 = xn3 & multm_reduce_sb148;
  assign multm_reduce_mulsc_mulb_cq149 = xn3 & multm_reduce_sb149;
  assign multm_reduce_mulsc_mulb_cq150 = xn3 & multm_reduce_sb150;
  assign multm_reduce_mulsc_mulb_cq151 = xn3 & multm_reduce_sb151;
  assign multm_reduce_mulsc_mulb_cq152 = xn3 & multm_reduce_sb152;
  assign multm_reduce_mulsc_mulb_cq153 = xn3 & multm_reduce_sb153;
  assign multm_reduce_mulsc_mulb_cq154 = xn3 & multm_reduce_sb154;
  assign multm_reduce_mulsc_mulb_cq155 = xn3 & multm_reduce_sb155;
  assign multm_reduce_mulsc_mulb_cq156 = xn3 & multm_reduce_sb156;
  assign multm_reduce_mulsc_mulb_cq157 = xn3 & multm_reduce_sb157;
  assign multm_reduce_mulsc_mulb_cq158 = xn3 & multm_reduce_sb158;
  assign multm_reduce_mulsc_mulb_cq159 = xn3 & multm_reduce_sb159;
  assign multm_reduce_mulsc_mulb_cq160 = xn3 & multm_reduce_sb160;
  assign multm_reduce_mulsc_mulb_cq161 = xn3 & multm_reduce_sb161;
  assign multm_reduce_mulsc_mulb_cq162 = xn3 & multm_reduce_sb162;
  assign multm_reduce_mulsc_mulb_cq163 = xn3 & multm_reduce_sb163;
  assign multm_reduce_mulsc_mulb_cq164 = xn3 & multm_reduce_sb164;
  assign multm_reduce_mulsc_mulb_cq165 = xn3 & multm_reduce_sb165;
  assign multm_reduce_mulsc_mulb_cq166 = xn3 & multm_reduce_sb166;
  assign multm_reduce_mulsc_mulb_cq167 = xn3 & multm_reduce_sb167;
  assign multm_reduce_mulsc_mulb_cq168 = xn3 & multm_reduce_sb168;
  assign multm_reduce_mulsc_mulb_cq169 = xn3 & multm_reduce_sb169;
  assign multm_reduce_mulsc_mulb_cq170 = xn3 & multm_reduce_sb170;
  assign multm_reduce_mulsc_mulb_cq171 = xn3 & multm_reduce_sb171;
  assign multm_reduce_mulsc_mulb_cq172 = xn3 & multm_reduce_sb172;
  assign multm_reduce_mulsc_mulb_cq173 = xn3 & multm_reduce_sb173;
  assign multm_reduce_mulsc_mulb_cq174 = xn3 & multm_reduce_sb174;
  assign multm_reduce_mulsc_mulb_cq175 = xn3 & multm_reduce_mulsc_mulb_cp175;
  assign multm_reduce_mulsc_mulb_cq176 = xn3 & multm_reduce_mulsc_mulb_cp176;
  assign multm_reduce_mulsc_mulb_cq177 = xn3 & multm_reduce_mulsc_mulb_cp177;
  assign multm_reduce_mulsc_mulb_cq178 = xn3 & multm_reduce_mulsc_mulb_cp178;
  assign multm_reduce_mulsc_mulb_cq179 = xn3 & multm_reduce_mulsc_mulb_cp179;
  assign multm_reduce_mulsc_mulb_cq180 = xn3 & multm_reduce_mulsc_mulb_cp180;
  assign multm_reduce_mulsc_mulb_cq181 = xn3 & multm_reduce_mulsc_mulb_cp181;
  assign multm_reduce_mulsc_mulb_cq182 = xn3 & multm_reduce_mulsc_mulb_cp182;
  assign multm_reduce_mulsc_mulb_cq183 = xn3 & multm_reduce_mulsc_mulb_cp183;
  assign multm_reduce_mulsc_mulb_pc0 = multm_reduce_mulsc_mulb_sq0 & multm_reduce_mulsc_mulb_yos0;
  assign multm_reduce_mulsc_mulb_pc1 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx0 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy0;
  assign multm_reduce_mulsc_mulb_pc2 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx1 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy1;
  assign multm_reduce_mulsc_mulb_pc3 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx2 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy2;
  assign multm_reduce_mulsc_mulb_pc4 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx3 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy3;
  assign multm_reduce_mulsc_mulb_pc5 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx4 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy4;
  assign multm_reduce_mulsc_mulb_pc6 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx5 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy5;
  assign multm_reduce_mulsc_mulb_pc7 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx6 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy6;
  assign multm_reduce_mulsc_mulb_pc8 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx7 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy7;
  assign multm_reduce_mulsc_mulb_pc9 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx8 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy8;
  assign multm_reduce_mulsc_mulb_pc10 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx9 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy9;
  assign multm_reduce_mulsc_mulb_pc11 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx10 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy10;
  assign multm_reduce_mulsc_mulb_pc12 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx11 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy11;
  assign multm_reduce_mulsc_mulb_pc13 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx12 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy12;
  assign multm_reduce_mulsc_mulb_pc14 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx13 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy13;
  assign multm_reduce_mulsc_mulb_pc15 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx14 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy14;
  assign multm_reduce_mulsc_mulb_pc16 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx15 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy15;
  assign multm_reduce_mulsc_mulb_pc17 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx16 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy16;
  assign multm_reduce_mulsc_mulb_pc18 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx17 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy17;
  assign multm_reduce_mulsc_mulb_pc19 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx18 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy18;
  assign multm_reduce_mulsc_mulb_pc20 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx19 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy19;
  assign multm_reduce_mulsc_mulb_pc21 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx20 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy20;
  assign multm_reduce_mulsc_mulb_pc22 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx21 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy21;
  assign multm_reduce_mulsc_mulb_pc23 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx22 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy22;
  assign multm_reduce_mulsc_mulb_pc24 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx23 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy23;
  assign multm_reduce_mulsc_mulb_pc25 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx24 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy24;
  assign multm_reduce_mulsc_mulb_pc26 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx25 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy25;
  assign multm_reduce_mulsc_mulb_pc27 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx26 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy26;
  assign multm_reduce_mulsc_mulb_pc28 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx27 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy27;
  assign multm_reduce_mulsc_mulb_pc29 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx28 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy28;
  assign multm_reduce_mulsc_mulb_pc30 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx29 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy29;
  assign multm_reduce_mulsc_mulb_pc31 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx30 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy30;
  assign multm_reduce_mulsc_mulb_pc32 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx31 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy31;
  assign multm_reduce_mulsc_mulb_pc33 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx32 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy32;
  assign multm_reduce_mulsc_mulb_pc34 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx33 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy33;
  assign multm_reduce_mulsc_mulb_pc35 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx34 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy34;
  assign multm_reduce_mulsc_mulb_pc36 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx35 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy35;
  assign multm_reduce_mulsc_mulb_pc37 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx36 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy36;
  assign multm_reduce_mulsc_mulb_pc38 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx37 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy37;
  assign multm_reduce_mulsc_mulb_pc39 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx38 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy38;
  assign multm_reduce_mulsc_mulb_pc40 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx39 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy39;
  assign multm_reduce_mulsc_mulb_pc41 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx40 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy40;
  assign multm_reduce_mulsc_mulb_pc42 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx41 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy41;
  assign multm_reduce_mulsc_mulb_pc43 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx42 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy42;
  assign multm_reduce_mulsc_mulb_pc44 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx43 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy43;
  assign multm_reduce_mulsc_mulb_pc45 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx44 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy44;
  assign multm_reduce_mulsc_mulb_pc46 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx45 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy45;
  assign multm_reduce_mulsc_mulb_pc47 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx46 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy46;
  assign multm_reduce_mulsc_mulb_pc48 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx47 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy47;
  assign multm_reduce_mulsc_mulb_pc49 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx48 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy48;
  assign multm_reduce_mulsc_mulb_pc50 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx49 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy49;
  assign multm_reduce_mulsc_mulb_pc51 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx50 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy50;
  assign multm_reduce_mulsc_mulb_pc52 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx51 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy51;
  assign multm_reduce_mulsc_mulb_pc53 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx52 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy52;
  assign multm_reduce_mulsc_mulb_pc54 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx53 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy53;
  assign multm_reduce_mulsc_mulb_pc55 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx54 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy54;
  assign multm_reduce_mulsc_mulb_pc56 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx55 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy55;
  assign multm_reduce_mulsc_mulb_pc57 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx56 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy56;
  assign multm_reduce_mulsc_mulb_pc58 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx57 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy57;
  assign multm_reduce_mulsc_mulb_pc59 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx58 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy58;
  assign multm_reduce_mulsc_mulb_pc60 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx59 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy59;
  assign multm_reduce_mulsc_mulb_pc61 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx60 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy60;
  assign multm_reduce_mulsc_mulb_pc62 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx61 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy61;
  assign multm_reduce_mulsc_mulb_pc63 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx62 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy62;
  assign multm_reduce_mulsc_mulb_pc64 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx63 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy63;
  assign multm_reduce_mulsc_mulb_pc65 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx64 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy64;
  assign multm_reduce_mulsc_mulb_pc66 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx65 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy65;
  assign multm_reduce_mulsc_mulb_pc67 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx66 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy66;
  assign multm_reduce_mulsc_mulb_pc68 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx67 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy67;
  assign multm_reduce_mulsc_mulb_pc69 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx68 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy68;
  assign multm_reduce_mulsc_mulb_pc70 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx69 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy69;
  assign multm_reduce_mulsc_mulb_pc71 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx70 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy70;
  assign multm_reduce_mulsc_mulb_pc72 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx71 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy71;
  assign multm_reduce_mulsc_mulb_pc73 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx72 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy72;
  assign multm_reduce_mulsc_mulb_pc74 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx73 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy73;
  assign multm_reduce_mulsc_mulb_pc75 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx74 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy74;
  assign multm_reduce_mulsc_mulb_pc76 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx75 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy75;
  assign multm_reduce_mulsc_mulb_pc77 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx76 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy76;
  assign multm_reduce_mulsc_mulb_pc78 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx77 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy77;
  assign multm_reduce_mulsc_mulb_pc79 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx78 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy78;
  assign multm_reduce_mulsc_mulb_pc80 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx79 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy79;
  assign multm_reduce_mulsc_mulb_pc81 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx80 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy80;
  assign multm_reduce_mulsc_mulb_pc82 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx81 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy81;
  assign multm_reduce_mulsc_mulb_pc83 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx82 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy82;
  assign multm_reduce_mulsc_mulb_pc84 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx83 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy83;
  assign multm_reduce_mulsc_mulb_pc85 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx84 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy84;
  assign multm_reduce_mulsc_mulb_pc86 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx85 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy85;
  assign multm_reduce_mulsc_mulb_pc87 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx86 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy86;
  assign multm_reduce_mulsc_mulb_pc88 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx87 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy87;
  assign multm_reduce_mulsc_mulb_pc89 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx88 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy88;
  assign multm_reduce_mulsc_mulb_pc90 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx89 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy89;
  assign multm_reduce_mulsc_mulb_pc91 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx90 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy90;
  assign multm_reduce_mulsc_mulb_pc92 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx91 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy91;
  assign multm_reduce_mulsc_mulb_pc93 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx92 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy92;
  assign multm_reduce_mulsc_mulb_pc94 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx93 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy93;
  assign multm_reduce_mulsc_mulb_pc95 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx94 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy94;
  assign multm_reduce_mulsc_mulb_pc96 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx95 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy95;
  assign multm_reduce_mulsc_mulb_pc97 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx96 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy96;
  assign multm_reduce_mulsc_mulb_pc98 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx97 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy97;
  assign multm_reduce_mulsc_mulb_pc99 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx98 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy98;
  assign multm_reduce_mulsc_mulb_pc100 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx99 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy99;
  assign multm_reduce_mulsc_mulb_pc101 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx100 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy100;
  assign multm_reduce_mulsc_mulb_pc102 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx101 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy101;
  assign multm_reduce_mulsc_mulb_pc103 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx102 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy102;
  assign multm_reduce_mulsc_mulb_pc104 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx103 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy103;
  assign multm_reduce_mulsc_mulb_pc105 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx104 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy104;
  assign multm_reduce_mulsc_mulb_pc106 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx105 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy105;
  assign multm_reduce_mulsc_mulb_pc107 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx106 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy106;
  assign multm_reduce_mulsc_mulb_pc108 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx107 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy107;
  assign multm_reduce_mulsc_mulb_pc109 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx108 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy108;
  assign multm_reduce_mulsc_mulb_pc110 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx109 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy109;
  assign multm_reduce_mulsc_mulb_pc111 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx110 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy110;
  assign multm_reduce_mulsc_mulb_pc112 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx111 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy111;
  assign multm_reduce_mulsc_mulb_pc113 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx112 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy112;
  assign multm_reduce_mulsc_mulb_pc114 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx113 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy113;
  assign multm_reduce_mulsc_mulb_pc115 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx114 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy114;
  assign multm_reduce_mulsc_mulb_pc116 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx115 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy115;
  assign multm_reduce_mulsc_mulb_pc117 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx116 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy116;
  assign multm_reduce_mulsc_mulb_pc118 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx117 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy117;
  assign multm_reduce_mulsc_mulb_pc119 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx118 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy118;
  assign multm_reduce_mulsc_mulb_pc120 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx119 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy119;
  assign multm_reduce_mulsc_mulb_pc121 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx120 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy120;
  assign multm_reduce_mulsc_mulb_pc122 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx121 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy121;
  assign multm_reduce_mulsc_mulb_pc123 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx122 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy122;
  assign multm_reduce_mulsc_mulb_pc124 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx123 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy123;
  assign multm_reduce_mulsc_mulb_pc125 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx124 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy124;
  assign multm_reduce_mulsc_mulb_pc126 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx125 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy125;
  assign multm_reduce_mulsc_mulb_pc127 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx126 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy126;
  assign multm_reduce_mulsc_mulb_pc128 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx127 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy127;
  assign multm_reduce_mulsc_mulb_pc129 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx128 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy128;
  assign multm_reduce_mulsc_mulb_pc130 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx129 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy129;
  assign multm_reduce_mulsc_mulb_pc131 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx130 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy130;
  assign multm_reduce_mulsc_mulb_pc132 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx131 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy131;
  assign multm_reduce_mulsc_mulb_pc133 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx132 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy132;
  assign multm_reduce_mulsc_mulb_pc134 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx133 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy133;
  assign multm_reduce_mulsc_mulb_pc135 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx134 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy134;
  assign multm_reduce_mulsc_mulb_pc136 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx135 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy135;
  assign multm_reduce_mulsc_mulb_pc137 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx136 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy136;
  assign multm_reduce_mulsc_mulb_pc138 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx137 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy137;
  assign multm_reduce_mulsc_mulb_pc139 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx138 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy138;
  assign multm_reduce_mulsc_mulb_pc140 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx139 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy139;
  assign multm_reduce_mulsc_mulb_pc141 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx140 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy140;
  assign multm_reduce_mulsc_mulb_pc142 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx141 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy141;
  assign multm_reduce_mulsc_mulb_pc143 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx142 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy142;
  assign multm_reduce_mulsc_mulb_pc144 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx143 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy143;
  assign multm_reduce_mulsc_mulb_pc145 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx144 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy144;
  assign multm_reduce_mulsc_mulb_pc146 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx145 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy145;
  assign multm_reduce_mulsc_mulb_pc147 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx146 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy146;
  assign multm_reduce_mulsc_mulb_pc148 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx147 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy147;
  assign multm_reduce_mulsc_mulb_pc149 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx148 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy148;
  assign multm_reduce_mulsc_mulb_pc150 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx149 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy149;
  assign multm_reduce_mulsc_mulb_pc151 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx150 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy150;
  assign multm_reduce_mulsc_mulb_pc152 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx151 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy151;
  assign multm_reduce_mulsc_mulb_pc153 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx152 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy152;
  assign multm_reduce_mulsc_mulb_pc154 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx153 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy153;
  assign multm_reduce_mulsc_mulb_pc155 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx154 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy154;
  assign multm_reduce_mulsc_mulb_pc156 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx155 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy155;
  assign multm_reduce_mulsc_mulb_pc157 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx156 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy156;
  assign multm_reduce_mulsc_mulb_pc158 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx157 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy157;
  assign multm_reduce_mulsc_mulb_pc159 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx158 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy158;
  assign multm_reduce_mulsc_mulb_pc160 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx159 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy159;
  assign multm_reduce_mulsc_mulb_pc161 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx160 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy160;
  assign multm_reduce_mulsc_mulb_pc162 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx161 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy161;
  assign multm_reduce_mulsc_mulb_pc163 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx162 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy162;
  assign multm_reduce_mulsc_mulb_pc164 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx163 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy163;
  assign multm_reduce_mulsc_mulb_pc165 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx164 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy164;
  assign multm_reduce_mulsc_mulb_pc166 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx165 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy165;
  assign multm_reduce_mulsc_mulb_pc167 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx166 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy166;
  assign multm_reduce_mulsc_mulb_pc168 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx167 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy167;
  assign multm_reduce_mulsc_mulb_pc169 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx168 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy168;
  assign multm_reduce_mulsc_mulb_pc170 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx169 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy169;
  assign multm_reduce_mulsc_mulb_pc171 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx170 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy170;
  assign multm_reduce_mulsc_mulb_pc172 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx171 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy171;
  assign multm_reduce_mulsc_mulb_pc173 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx172 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy172;
  assign multm_reduce_mulsc_mulb_pc174 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx173 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy173;
  assign multm_reduce_mulsc_mulb_pc175 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx174 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy174;
  assign multm_reduce_mulsc_mulb_pc176 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx175 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy175;
  assign multm_reduce_mulsc_mulb_pc177 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx176 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy176;
  assign multm_reduce_mulsc_mulb_pc178 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx177 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy177;
  assign multm_reduce_mulsc_mulb_pc179 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx178 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy178;
  assign multm_reduce_mulsc_mulb_pc180 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx179 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy179;
  assign multm_reduce_mulsc_mulb_pc181 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx180 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy180;
  assign multm_reduce_mulsc_mulb_pc182 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx181 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy181;
  assign multm_reduce_mulsc_mulb_pc183 = multm_reduce_mulsc_mulb_add3b0_maj3b_or3b_wx182 | multm_reduce_mulsc_mulb_add3b0_maj3b_xy182;
  assign multm_reduce_mulsc_mulb_ps0 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx0 ^ multm_reduce_mulsc_mulb_yos1;
  assign multm_reduce_mulsc_mulb_ps1 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx1 ^ multm_reduce_mulsc_mulb_yos2;
  assign multm_reduce_mulsc_mulb_ps2 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx2 ^ multm_reduce_mulsc_mulb_yos3;
  assign multm_reduce_mulsc_mulb_ps3 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx3 ^ multm_reduce_mulsc_mulb_yos4;
  assign multm_reduce_mulsc_mulb_ps4 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx4 ^ multm_reduce_mulsc_mulb_yos5;
  assign multm_reduce_mulsc_mulb_ps5 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx5 ^ multm_reduce_mulsc_mulb_yos6;
  assign multm_reduce_mulsc_mulb_ps6 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx6 ^ multm_reduce_mulsc_mulb_yos7;
  assign multm_reduce_mulsc_mulb_ps7 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx7 ^ multm_reduce_mulsc_mulb_yos8;
  assign multm_reduce_mulsc_mulb_ps8 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx8 ^ multm_reduce_mulsc_mulb_yos9;
  assign multm_reduce_mulsc_mulb_ps9 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx9 ^ multm_reduce_mulsc_mulb_yos10;
  assign multm_reduce_mulsc_mulb_ps10 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx10 ^ multm_reduce_mulsc_mulb_yos11;
  assign multm_reduce_mulsc_mulb_ps11 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx11 ^ multm_reduce_mulsc_mulb_yos12;
  assign multm_reduce_mulsc_mulb_ps12 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx12 ^ multm_reduce_mulsc_mulb_yos13;
  assign multm_reduce_mulsc_mulb_ps13 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx13 ^ multm_reduce_mulsc_mulb_yos14;
  assign multm_reduce_mulsc_mulb_ps14 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx14 ^ multm_reduce_mulsc_mulb_yos15;
  assign multm_reduce_mulsc_mulb_ps15 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx15 ^ multm_reduce_mulsc_mulb_yos16;
  assign multm_reduce_mulsc_mulb_ps16 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx16 ^ multm_reduce_mulsc_mulb_yos17;
  assign multm_reduce_mulsc_mulb_ps17 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx17 ^ multm_reduce_mulsc_mulb_yos18;
  assign multm_reduce_mulsc_mulb_ps18 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx18 ^ multm_reduce_mulsc_mulb_yos19;
  assign multm_reduce_mulsc_mulb_ps19 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx19 ^ multm_reduce_mulsc_mulb_yos20;
  assign multm_reduce_mulsc_mulb_ps20 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx20 ^ multm_reduce_mulsc_mulb_yos21;
  assign multm_reduce_mulsc_mulb_ps21 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx21 ^ multm_reduce_mulsc_mulb_yos22;
  assign multm_reduce_mulsc_mulb_ps22 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx22 ^ multm_reduce_mulsc_mulb_yos23;
  assign multm_reduce_mulsc_mulb_ps23 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx23 ^ multm_reduce_mulsc_mulb_yos24;
  assign multm_reduce_mulsc_mulb_ps24 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx24 ^ multm_reduce_mulsc_mulb_yos25;
  assign multm_reduce_mulsc_mulb_ps25 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx25 ^ multm_reduce_mulsc_mulb_yos26;
  assign multm_reduce_mulsc_mulb_ps26 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx26 ^ multm_reduce_mulsc_mulb_yos27;
  assign multm_reduce_mulsc_mulb_ps27 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx27 ^ multm_reduce_mulsc_mulb_yos28;
  assign multm_reduce_mulsc_mulb_ps28 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx28 ^ multm_reduce_mulsc_mulb_yos29;
  assign multm_reduce_mulsc_mulb_ps29 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx29 ^ multm_reduce_mulsc_mulb_yos30;
  assign multm_reduce_mulsc_mulb_ps30 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx30 ^ multm_reduce_mulsc_mulb_yos31;
  assign multm_reduce_mulsc_mulb_ps31 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx31 ^ multm_reduce_mulsc_mulb_yos32;
  assign multm_reduce_mulsc_mulb_ps32 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx32 ^ multm_reduce_mulsc_mulb_yos33;
  assign multm_reduce_mulsc_mulb_ps33 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx33 ^ multm_reduce_mulsc_mulb_yos34;
  assign multm_reduce_mulsc_mulb_ps34 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx34 ^ multm_reduce_mulsc_mulb_yos35;
  assign multm_reduce_mulsc_mulb_ps35 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx35 ^ multm_reduce_mulsc_mulb_yos36;
  assign multm_reduce_mulsc_mulb_ps36 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx36 ^ multm_reduce_mulsc_mulb_yos37;
  assign multm_reduce_mulsc_mulb_ps37 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx37 ^ multm_reduce_mulsc_mulb_yos38;
  assign multm_reduce_mulsc_mulb_ps38 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx38 ^ multm_reduce_mulsc_mulb_yos39;
  assign multm_reduce_mulsc_mulb_ps39 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx39 ^ multm_reduce_mulsc_mulb_yos40;
  assign multm_reduce_mulsc_mulb_ps40 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx40 ^ multm_reduce_mulsc_mulb_yos41;
  assign multm_reduce_mulsc_mulb_ps41 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx41 ^ multm_reduce_mulsc_mulb_yos42;
  assign multm_reduce_mulsc_mulb_ps42 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx42 ^ multm_reduce_mulsc_mulb_yos43;
  assign multm_reduce_mulsc_mulb_ps43 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx43 ^ multm_reduce_mulsc_mulb_yos44;
  assign multm_reduce_mulsc_mulb_ps44 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx44 ^ multm_reduce_mulsc_mulb_yos45;
  assign multm_reduce_mulsc_mulb_ps45 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx45 ^ multm_reduce_mulsc_mulb_yos46;
  assign multm_reduce_mulsc_mulb_ps46 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx46 ^ multm_reduce_mulsc_mulb_yos47;
  assign multm_reduce_mulsc_mulb_ps47 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx47 ^ multm_reduce_mulsc_mulb_yos48;
  assign multm_reduce_mulsc_mulb_ps48 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx48 ^ multm_reduce_mulsc_mulb_yos49;
  assign multm_reduce_mulsc_mulb_ps49 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx49 ^ multm_reduce_mulsc_mulb_yos50;
  assign multm_reduce_mulsc_mulb_ps50 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx50 ^ multm_reduce_mulsc_mulb_yos51;
  assign multm_reduce_mulsc_mulb_ps51 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx51 ^ multm_reduce_mulsc_mulb_yos52;
  assign multm_reduce_mulsc_mulb_ps52 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx52 ^ multm_reduce_mulsc_mulb_yos53;
  assign multm_reduce_mulsc_mulb_ps53 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx53 ^ multm_reduce_mulsc_mulb_yos54;
  assign multm_reduce_mulsc_mulb_ps54 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx54 ^ multm_reduce_mulsc_mulb_yos55;
  assign multm_reduce_mulsc_mulb_ps55 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx55 ^ multm_reduce_mulsc_mulb_yos56;
  assign multm_reduce_mulsc_mulb_ps56 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx56 ^ multm_reduce_mulsc_mulb_yos57;
  assign multm_reduce_mulsc_mulb_ps57 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx57 ^ multm_reduce_mulsc_mulb_yos58;
  assign multm_reduce_mulsc_mulb_ps58 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx58 ^ multm_reduce_mulsc_mulb_yos59;
  assign multm_reduce_mulsc_mulb_ps59 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx59 ^ multm_reduce_mulsc_mulb_yos60;
  assign multm_reduce_mulsc_mulb_ps60 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx60 ^ multm_reduce_mulsc_mulb_yos61;
  assign multm_reduce_mulsc_mulb_ps61 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx61 ^ multm_reduce_mulsc_mulb_yos62;
  assign multm_reduce_mulsc_mulb_ps62 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx62 ^ multm_reduce_mulsc_mulb_yos63;
  assign multm_reduce_mulsc_mulb_ps63 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx63 ^ multm_reduce_mulsc_mulb_yos64;
  assign multm_reduce_mulsc_mulb_ps64 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx64 ^ multm_reduce_mulsc_mulb_yos65;
  assign multm_reduce_mulsc_mulb_ps65 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx65 ^ multm_reduce_mulsc_mulb_yos66;
  assign multm_reduce_mulsc_mulb_ps66 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx66 ^ multm_reduce_mulsc_mulb_yos67;
  assign multm_reduce_mulsc_mulb_ps67 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx67 ^ multm_reduce_mulsc_mulb_yos68;
  assign multm_reduce_mulsc_mulb_ps68 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx68 ^ multm_reduce_mulsc_mulb_yos69;
  assign multm_reduce_mulsc_mulb_ps69 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx69 ^ multm_reduce_mulsc_mulb_yos70;
  assign multm_reduce_mulsc_mulb_ps70 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx70 ^ multm_reduce_mulsc_mulb_yos71;
  assign multm_reduce_mulsc_mulb_ps71 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx71 ^ multm_reduce_mulsc_mulb_yos72;
  assign multm_reduce_mulsc_mulb_ps72 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx72 ^ multm_reduce_mulsc_mulb_yos73;
  assign multm_reduce_mulsc_mulb_ps73 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx73 ^ multm_reduce_mulsc_mulb_yos74;
  assign multm_reduce_mulsc_mulb_ps74 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx74 ^ multm_reduce_mulsc_mulb_yos75;
  assign multm_reduce_mulsc_mulb_ps75 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx75 ^ multm_reduce_mulsc_mulb_yos76;
  assign multm_reduce_mulsc_mulb_ps76 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx76 ^ multm_reduce_mulsc_mulb_yos77;
  assign multm_reduce_mulsc_mulb_ps77 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx77 ^ multm_reduce_mulsc_mulb_yos78;
  assign multm_reduce_mulsc_mulb_ps78 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx78 ^ multm_reduce_mulsc_mulb_yos79;
  assign multm_reduce_mulsc_mulb_ps79 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx79 ^ multm_reduce_mulsc_mulb_yos80;
  assign multm_reduce_mulsc_mulb_ps80 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx80 ^ multm_reduce_mulsc_mulb_yos81;
  assign multm_reduce_mulsc_mulb_ps81 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx81 ^ multm_reduce_mulsc_mulb_yos82;
  assign multm_reduce_mulsc_mulb_ps82 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx82 ^ multm_reduce_mulsc_mulb_yos83;
  assign multm_reduce_mulsc_mulb_ps83 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx83 ^ multm_reduce_mulsc_mulb_yos84;
  assign multm_reduce_mulsc_mulb_ps84 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx84 ^ multm_reduce_mulsc_mulb_yos85;
  assign multm_reduce_mulsc_mulb_ps85 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx85 ^ multm_reduce_mulsc_mulb_yos86;
  assign multm_reduce_mulsc_mulb_ps86 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx86 ^ multm_reduce_mulsc_mulb_yos87;
  assign multm_reduce_mulsc_mulb_ps87 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx87 ^ multm_reduce_mulsc_mulb_yos88;
  assign multm_reduce_mulsc_mulb_ps88 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx88 ^ multm_reduce_mulsc_mulb_yos89;
  assign multm_reduce_mulsc_mulb_ps89 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx89 ^ multm_reduce_mulsc_mulb_yos90;
  assign multm_reduce_mulsc_mulb_ps90 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx90 ^ multm_reduce_mulsc_mulb_yos91;
  assign multm_reduce_mulsc_mulb_ps91 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx91 ^ multm_reduce_mulsc_mulb_yos92;
  assign multm_reduce_mulsc_mulb_ps92 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx92 ^ multm_reduce_mulsc_mulb_yos93;
  assign multm_reduce_mulsc_mulb_ps93 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx93 ^ multm_reduce_mulsc_mulb_yos94;
  assign multm_reduce_mulsc_mulb_ps94 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx94 ^ multm_reduce_mulsc_mulb_yos95;
  assign multm_reduce_mulsc_mulb_ps95 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx95 ^ multm_reduce_mulsc_mulb_yos96;
  assign multm_reduce_mulsc_mulb_ps96 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx96 ^ multm_reduce_mulsc_mulb_yos97;
  assign multm_reduce_mulsc_mulb_ps97 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx97 ^ multm_reduce_mulsc_mulb_yos98;
  assign multm_reduce_mulsc_mulb_ps98 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx98 ^ multm_reduce_mulsc_mulb_yos99;
  assign multm_reduce_mulsc_mulb_ps99 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx99 ^ multm_reduce_mulsc_mulb_yos100;
  assign multm_reduce_mulsc_mulb_ps100 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx100 ^ multm_reduce_mulsc_mulb_yos101;
  assign multm_reduce_mulsc_mulb_ps101 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx101 ^ multm_reduce_mulsc_mulb_yos102;
  assign multm_reduce_mulsc_mulb_ps102 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx102 ^ multm_reduce_mulsc_mulb_yos103;
  assign multm_reduce_mulsc_mulb_ps103 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx103 ^ multm_reduce_mulsc_mulb_yos104;
  assign multm_reduce_mulsc_mulb_ps104 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx104 ^ multm_reduce_mulsc_mulb_yos105;
  assign multm_reduce_mulsc_mulb_ps105 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx105 ^ multm_reduce_mulsc_mulb_yos106;
  assign multm_reduce_mulsc_mulb_ps106 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx106 ^ multm_reduce_mulsc_mulb_yos107;
  assign multm_reduce_mulsc_mulb_ps107 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx107 ^ multm_reduce_mulsc_mulb_yos108;
  assign multm_reduce_mulsc_mulb_ps108 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx108 ^ multm_reduce_mulsc_mulb_yos109;
  assign multm_reduce_mulsc_mulb_ps109 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx109 ^ multm_reduce_mulsc_mulb_yos110;
  assign multm_reduce_mulsc_mulb_ps110 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx110 ^ multm_reduce_mulsc_mulb_yos111;
  assign multm_reduce_mulsc_mulb_ps111 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx111 ^ multm_reduce_mulsc_mulb_yos112;
  assign multm_reduce_mulsc_mulb_ps112 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx112 ^ multm_reduce_mulsc_mulb_yos113;
  assign multm_reduce_mulsc_mulb_ps113 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx113 ^ multm_reduce_mulsc_mulb_yos114;
  assign multm_reduce_mulsc_mulb_ps114 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx114 ^ multm_reduce_mulsc_mulb_yos115;
  assign multm_reduce_mulsc_mulb_ps115 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx115 ^ multm_reduce_mulsc_mulb_yos116;
  assign multm_reduce_mulsc_mulb_ps116 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx116 ^ multm_reduce_mulsc_mulb_yos117;
  assign multm_reduce_mulsc_mulb_ps117 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx117 ^ multm_reduce_mulsc_mulb_yos118;
  assign multm_reduce_mulsc_mulb_ps118 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx118 ^ multm_reduce_mulsc_mulb_yos119;
  assign multm_reduce_mulsc_mulb_ps119 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx119 ^ multm_reduce_mulsc_mulb_yos120;
  assign multm_reduce_mulsc_mulb_ps120 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx120 ^ multm_reduce_mulsc_mulb_yos121;
  assign multm_reduce_mulsc_mulb_ps121 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx121 ^ multm_reduce_mulsc_mulb_yos122;
  assign multm_reduce_mulsc_mulb_ps122 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx122 ^ multm_reduce_mulsc_mulb_yos123;
  assign multm_reduce_mulsc_mulb_ps123 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx123 ^ multm_reduce_mulsc_mulb_yos124;
  assign multm_reduce_mulsc_mulb_ps124 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx124 ^ multm_reduce_mulsc_mulb_yos125;
  assign multm_reduce_mulsc_mulb_ps125 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx125 ^ multm_reduce_mulsc_mulb_yos126;
  assign multm_reduce_mulsc_mulb_ps126 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx126 ^ multm_reduce_mulsc_mulb_yos127;
  assign multm_reduce_mulsc_mulb_ps127 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx127 ^ multm_reduce_mulsc_mulb_yos128;
  assign multm_reduce_mulsc_mulb_ps128 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx128 ^ multm_reduce_mulsc_mulb_yos129;
  assign multm_reduce_mulsc_mulb_ps129 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx129 ^ multm_reduce_mulsc_mulb_yos130;
  assign multm_reduce_mulsc_mulb_ps130 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx130 ^ multm_reduce_mulsc_mulb_yos131;
  assign multm_reduce_mulsc_mulb_ps131 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx131 ^ multm_reduce_mulsc_mulb_yos132;
  assign multm_reduce_mulsc_mulb_ps132 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx132 ^ multm_reduce_mulsc_mulb_yos133;
  assign multm_reduce_mulsc_mulb_ps133 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx133 ^ multm_reduce_mulsc_mulb_yos134;
  assign multm_reduce_mulsc_mulb_ps134 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx134 ^ multm_reduce_mulsc_mulb_yos135;
  assign multm_reduce_mulsc_mulb_ps135 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx135 ^ multm_reduce_mulsc_mulb_yos136;
  assign multm_reduce_mulsc_mulb_ps136 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx136 ^ multm_reduce_mulsc_mulb_yos137;
  assign multm_reduce_mulsc_mulb_ps137 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx137 ^ multm_reduce_mulsc_mulb_yos138;
  assign multm_reduce_mulsc_mulb_ps138 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx138 ^ multm_reduce_mulsc_mulb_yos139;
  assign multm_reduce_mulsc_mulb_ps139 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx139 ^ multm_reduce_mulsc_mulb_yos140;
  assign multm_reduce_mulsc_mulb_ps140 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx140 ^ multm_reduce_mulsc_mulb_yos141;
  assign multm_reduce_mulsc_mulb_ps141 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx141 ^ multm_reduce_mulsc_mulb_yos142;
  assign multm_reduce_mulsc_mulb_ps142 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx142 ^ multm_reduce_mulsc_mulb_yos143;
  assign multm_reduce_mulsc_mulb_ps143 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx143 ^ multm_reduce_mulsc_mulb_yos144;
  assign multm_reduce_mulsc_mulb_ps144 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx144 ^ multm_reduce_mulsc_mulb_yos145;
  assign multm_reduce_mulsc_mulb_ps145 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx145 ^ multm_reduce_mulsc_mulb_yos146;
  assign multm_reduce_mulsc_mulb_ps146 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx146 ^ multm_reduce_mulsc_mulb_yos147;
  assign multm_reduce_mulsc_mulb_ps147 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx147 ^ multm_reduce_mulsc_mulb_yos148;
  assign multm_reduce_mulsc_mulb_ps148 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx148 ^ multm_reduce_mulsc_mulb_yos149;
  assign multm_reduce_mulsc_mulb_ps149 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx149 ^ multm_reduce_mulsc_mulb_yos150;
  assign multm_reduce_mulsc_mulb_ps150 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx150 ^ multm_reduce_mulsc_mulb_yos151;
  assign multm_reduce_mulsc_mulb_ps151 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx151 ^ multm_reduce_mulsc_mulb_yos152;
  assign multm_reduce_mulsc_mulb_ps152 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx152 ^ multm_reduce_mulsc_mulb_yos153;
  assign multm_reduce_mulsc_mulb_ps153 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx153 ^ multm_reduce_mulsc_mulb_yos154;
  assign multm_reduce_mulsc_mulb_ps154 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx154 ^ multm_reduce_mulsc_mulb_yos155;
  assign multm_reduce_mulsc_mulb_ps155 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx155 ^ multm_reduce_mulsc_mulb_yos156;
  assign multm_reduce_mulsc_mulb_ps156 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx156 ^ multm_reduce_mulsc_mulb_yos157;
  assign multm_reduce_mulsc_mulb_ps157 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx157 ^ multm_reduce_mulsc_mulb_yos158;
  assign multm_reduce_mulsc_mulb_ps158 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx158 ^ multm_reduce_mulsc_mulb_yos159;
  assign multm_reduce_mulsc_mulb_ps159 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx159 ^ multm_reduce_mulsc_mulb_yos160;
  assign multm_reduce_mulsc_mulb_ps160 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx160 ^ multm_reduce_mulsc_mulb_yos161;
  assign multm_reduce_mulsc_mulb_ps161 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx161 ^ multm_reduce_mulsc_mulb_yos162;
  assign multm_reduce_mulsc_mulb_ps162 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx162 ^ multm_reduce_mulsc_mulb_yos163;
  assign multm_reduce_mulsc_mulb_ps163 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx163 ^ multm_reduce_mulsc_mulb_yos164;
  assign multm_reduce_mulsc_mulb_ps164 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx164 ^ multm_reduce_mulsc_mulb_yos165;
  assign multm_reduce_mulsc_mulb_ps165 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx165 ^ multm_reduce_mulsc_mulb_yos166;
  assign multm_reduce_mulsc_mulb_ps166 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx166 ^ multm_reduce_mulsc_mulb_yos167;
  assign multm_reduce_mulsc_mulb_ps167 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx167 ^ multm_reduce_mulsc_mulb_yos168;
  assign multm_reduce_mulsc_mulb_ps168 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx168 ^ multm_reduce_mulsc_mulb_yos169;
  assign multm_reduce_mulsc_mulb_ps169 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx169 ^ multm_reduce_mulsc_mulb_yos170;
  assign multm_reduce_mulsc_mulb_ps170 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx170 ^ multm_reduce_mulsc_mulb_yos171;
  assign multm_reduce_mulsc_mulb_ps171 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx171 ^ multm_reduce_mulsc_mulb_yos172;
  assign multm_reduce_mulsc_mulb_ps172 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx172 ^ multm_reduce_mulsc_mulb_yos173;
  assign multm_reduce_mulsc_mulb_ps173 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx173 ^ multm_reduce_mulsc_mulb_yos174;
  assign multm_reduce_mulsc_mulb_ps174 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx174 ^ multm_reduce_mulsc_mulb_yos175;
  assign multm_reduce_mulsc_mulb_ps175 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx175 ^ multm_reduce_mulsc_mulb_yos176;
  assign multm_reduce_mulsc_mulb_ps176 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx176 ^ multm_reduce_mulsc_mulb_yos177;
  assign multm_reduce_mulsc_mulb_ps177 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx177 ^ multm_reduce_mulsc_mulb_yos178;
  assign multm_reduce_mulsc_mulb_ps178 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx178 ^ multm_reduce_mulsc_mulb_yos179;
  assign multm_reduce_mulsc_mulb_ps179 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx179 ^ multm_reduce_mulsc_mulb_yos180;
  assign multm_reduce_mulsc_mulb_ps180 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx180 ^ multm_reduce_mulsc_mulb_yos181;
  assign multm_reduce_mulsc_mulb_ps181 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx181 ^ multm_reduce_mulsc_mulb_yos182;
  assign multm_reduce_mulsc_mulb_ps182 = multm_reduce_mulsc_mulb_add3b0_xor3b_wx182 ^ multm_reduce_mulsc_mulb_yos183;
  assign multm_reduce_mulsc_mulb_sq0 = xn3 & multm_reduce_sa10;
  assign multm_reduce_mulsc_mulb_sq1 = xn3 & multm_reduce_sa11;
  assign multm_reduce_mulsc_mulb_sq2 = xn3 & multm_reduce_sa12;
  assign multm_reduce_mulsc_mulb_sq3 = xn3 & multm_reduce_sa13;
  assign multm_reduce_mulsc_mulb_sq4 = xn3 & multm_reduce_sa14;
  assign multm_reduce_mulsc_mulb_sq5 = xn3 & multm_reduce_sa15;
  assign multm_reduce_mulsc_mulb_sq6 = xn3 & multm_reduce_sa16;
  assign multm_reduce_mulsc_mulb_sq7 = xn3 & multm_reduce_sa17;
  assign multm_reduce_mulsc_mulb_sq8 = xn3 & multm_reduce_sa18;
  assign multm_reduce_mulsc_mulb_sq9 = xn3 & multm_reduce_sa19;
  assign multm_reduce_mulsc_mulb_sq10 = xn3 & multm_reduce_sa20;
  assign multm_reduce_mulsc_mulb_sq11 = xn3 & multm_reduce_sa21;
  assign multm_reduce_mulsc_mulb_sq12 = xn3 & multm_reduce_sa22;
  assign multm_reduce_mulsc_mulb_sq13 = xn3 & multm_reduce_sa23;
  assign multm_reduce_mulsc_mulb_sq14 = xn3 & multm_reduce_sa24;
  assign multm_reduce_mulsc_mulb_sq15 = xn3 & multm_reduce_sa25;
  assign multm_reduce_mulsc_mulb_sq16 = xn3 & multm_reduce_sa26;
  assign multm_reduce_mulsc_mulb_sq17 = xn3 & multm_reduce_sa27;
  assign multm_reduce_mulsc_mulb_sq18 = xn3 & multm_reduce_sa28;
  assign multm_reduce_mulsc_mulb_sq19 = xn3 & multm_reduce_sa29;
  assign multm_reduce_mulsc_mulb_sq20 = xn3 & multm_reduce_sa30;
  assign multm_reduce_mulsc_mulb_sq21 = xn3 & multm_reduce_sa31;
  assign multm_reduce_mulsc_mulb_sq22 = xn3 & multm_reduce_sa32;
  assign multm_reduce_mulsc_mulb_sq23 = xn3 & multm_reduce_sa33;
  assign multm_reduce_mulsc_mulb_sq24 = xn3 & multm_reduce_sa34;
  assign multm_reduce_mulsc_mulb_sq25 = xn3 & multm_reduce_sa35;
  assign multm_reduce_mulsc_mulb_sq26 = xn3 & multm_reduce_sa36;
  assign multm_reduce_mulsc_mulb_sq27 = xn3 & multm_reduce_sa37;
  assign multm_reduce_mulsc_mulb_sq28 = xn3 & multm_reduce_sa38;
  assign multm_reduce_mulsc_mulb_sq29 = xn3 & multm_reduce_sa39;
  assign multm_reduce_mulsc_mulb_sq30 = xn3 & multm_reduce_sa40;
  assign multm_reduce_mulsc_mulb_sq31 = xn3 & multm_reduce_sa41;
  assign multm_reduce_mulsc_mulb_sq32 = xn3 & multm_reduce_sa42;
  assign multm_reduce_mulsc_mulb_sq33 = xn3 & multm_reduce_sa43;
  assign multm_reduce_mulsc_mulb_sq34 = xn3 & multm_reduce_sa44;
  assign multm_reduce_mulsc_mulb_sq35 = xn3 & multm_reduce_sa45;
  assign multm_reduce_mulsc_mulb_sq36 = xn3 & multm_reduce_sa46;
  assign multm_reduce_mulsc_mulb_sq37 = xn3 & multm_reduce_sa47;
  assign multm_reduce_mulsc_mulb_sq38 = xn3 & multm_reduce_sa48;
  assign multm_reduce_mulsc_mulb_sq39 = xn3 & multm_reduce_sa49;
  assign multm_reduce_mulsc_mulb_sq40 = xn3 & multm_reduce_sa50;
  assign multm_reduce_mulsc_mulb_sq41 = xn3 & multm_reduce_sa51;
  assign multm_reduce_mulsc_mulb_sq42 = xn3 & multm_reduce_sa52;
  assign multm_reduce_mulsc_mulb_sq43 = xn3 & multm_reduce_sa53;
  assign multm_reduce_mulsc_mulb_sq44 = xn3 & multm_reduce_sa54;
  assign multm_reduce_mulsc_mulb_sq45 = xn3 & multm_reduce_sa55;
  assign multm_reduce_mulsc_mulb_sq46 = xn3 & multm_reduce_sa56;
  assign multm_reduce_mulsc_mulb_sq47 = xn3 & multm_reduce_sa57;
  assign multm_reduce_mulsc_mulb_sq48 = xn3 & multm_reduce_sa58;
  assign multm_reduce_mulsc_mulb_sq49 = xn3 & multm_reduce_sa59;
  assign multm_reduce_mulsc_mulb_sq50 = xn3 & multm_reduce_sa60;
  assign multm_reduce_mulsc_mulb_sq51 = xn3 & multm_reduce_sa61;
  assign multm_reduce_mulsc_mulb_sq52 = xn3 & multm_reduce_sa62;
  assign multm_reduce_mulsc_mulb_sq53 = xn3 & multm_reduce_sa63;
  assign multm_reduce_mulsc_mulb_sq54 = xn3 & multm_reduce_sa64;
  assign multm_reduce_mulsc_mulb_sq55 = xn3 & multm_reduce_sa65;
  assign multm_reduce_mulsc_mulb_sq56 = xn3 & multm_reduce_sa66;
  assign multm_reduce_mulsc_mulb_sq57 = xn3 & multm_reduce_sa67;
  assign multm_reduce_mulsc_mulb_sq58 = xn3 & multm_reduce_sa68;
  assign multm_reduce_mulsc_mulb_sq59 = xn3 & multm_reduce_sa69;
  assign multm_reduce_mulsc_mulb_sq60 = xn3 & multm_reduce_sa70;
  assign multm_reduce_mulsc_mulb_sq61 = xn3 & multm_reduce_sa71;
  assign multm_reduce_mulsc_mulb_sq62 = xn3 & multm_reduce_sa72;
  assign multm_reduce_mulsc_mulb_sq63 = xn3 & multm_reduce_sa73;
  assign multm_reduce_mulsc_mulb_sq64 = xn3 & multm_reduce_sa74;
  assign multm_reduce_mulsc_mulb_sq65 = xn3 & multm_reduce_sa75;
  assign multm_reduce_mulsc_mulb_sq66 = xn3 & multm_reduce_sa76;
  assign multm_reduce_mulsc_mulb_sq67 = xn3 & multm_reduce_sa77;
  assign multm_reduce_mulsc_mulb_sq68 = xn3 & multm_reduce_sa78;
  assign multm_reduce_mulsc_mulb_sq69 = xn3 & multm_reduce_sa79;
  assign multm_reduce_mulsc_mulb_sq70 = xn3 & multm_reduce_sa80;
  assign multm_reduce_mulsc_mulb_sq71 = xn3 & multm_reduce_sa81;
  assign multm_reduce_mulsc_mulb_sq72 = xn3 & multm_reduce_sa82;
  assign multm_reduce_mulsc_mulb_sq73 = xn3 & multm_reduce_sa83;
  assign multm_reduce_mulsc_mulb_sq74 = xn3 & multm_reduce_sa84;
  assign multm_reduce_mulsc_mulb_sq75 = xn3 & multm_reduce_sa85;
  assign multm_reduce_mulsc_mulb_sq76 = xn3 & multm_reduce_sa86;
  assign multm_reduce_mulsc_mulb_sq77 = xn3 & multm_reduce_sa87;
  assign multm_reduce_mulsc_mulb_sq78 = xn3 & multm_reduce_sa88;
  assign multm_reduce_mulsc_mulb_sq79 = xn3 & multm_reduce_sa89;
  assign multm_reduce_mulsc_mulb_sq80 = xn3 & multm_reduce_sa90;
  assign multm_reduce_mulsc_mulb_sq81 = xn3 & multm_reduce_sa91;
  assign multm_reduce_mulsc_mulb_sq82 = xn3 & multm_reduce_sa92;
  assign multm_reduce_mulsc_mulb_sq83 = xn3 & multm_reduce_sa93;
  assign multm_reduce_mulsc_mulb_sq84 = xn3 & multm_reduce_sa94;
  assign multm_reduce_mulsc_mulb_sq85 = xn3 & multm_reduce_sa95;
  assign multm_reduce_mulsc_mulb_sq86 = xn3 & multm_reduce_sa96;
  assign multm_reduce_mulsc_mulb_sq87 = xn3 & multm_reduce_sa97;
  assign multm_reduce_mulsc_mulb_sq88 = xn3 & multm_reduce_sa98;
  assign multm_reduce_mulsc_mulb_sq89 = xn3 & multm_reduce_sa99;
  assign multm_reduce_mulsc_mulb_sq90 = xn3 & multm_reduce_sa100;
  assign multm_reduce_mulsc_mulb_sq91 = xn3 & multm_reduce_sa101;
  assign multm_reduce_mulsc_mulb_sq92 = xn3 & multm_reduce_sa102;
  assign multm_reduce_mulsc_mulb_sq93 = xn3 & multm_reduce_sa103;
  assign multm_reduce_mulsc_mulb_sq94 = xn3 & multm_reduce_sa104;
  assign multm_reduce_mulsc_mulb_sq95 = xn3 & multm_reduce_sa105;
  assign multm_reduce_mulsc_mulb_sq96 = xn3 & multm_reduce_sa106;
  assign multm_reduce_mulsc_mulb_sq97 = xn3 & multm_reduce_sa107;
  assign multm_reduce_mulsc_mulb_sq98 = xn3 & multm_reduce_sa108;
  assign multm_reduce_mulsc_mulb_sq99 = xn3 & multm_reduce_sa109;
  assign multm_reduce_mulsc_mulb_sq100 = xn3 & multm_reduce_sa110;
  assign multm_reduce_mulsc_mulb_sq101 = xn3 & multm_reduce_sa111;
  assign multm_reduce_mulsc_mulb_sq102 = xn3 & multm_reduce_sa112;
  assign multm_reduce_mulsc_mulb_sq103 = xn3 & multm_reduce_sa113;
  assign multm_reduce_mulsc_mulb_sq104 = xn3 & multm_reduce_sa114;
  assign multm_reduce_mulsc_mulb_sq105 = xn3 & multm_reduce_sa115;
  assign multm_reduce_mulsc_mulb_sq106 = xn3 & multm_reduce_sa116;
  assign multm_reduce_mulsc_mulb_sq107 = xn3 & multm_reduce_sa117;
  assign multm_reduce_mulsc_mulb_sq108 = xn3 & multm_reduce_sa118;
  assign multm_reduce_mulsc_mulb_sq109 = xn3 & multm_reduce_sa119;
  assign multm_reduce_mulsc_mulb_sq110 = xn3 & multm_reduce_sa120;
  assign multm_reduce_mulsc_mulb_sq111 = xn3 & multm_reduce_sa121;
  assign multm_reduce_mulsc_mulb_sq112 = xn3 & multm_reduce_sa122;
  assign multm_reduce_mulsc_mulb_sq113 = xn3 & multm_reduce_sa123;
  assign multm_reduce_mulsc_mulb_sq114 = xn3 & multm_reduce_sa124;
  assign multm_reduce_mulsc_mulb_sq115 = xn3 & multm_reduce_sa125;
  assign multm_reduce_mulsc_mulb_sq116 = xn3 & multm_reduce_sa126;
  assign multm_reduce_mulsc_mulb_sq117 = xn3 & multm_reduce_sa127;
  assign multm_reduce_mulsc_mulb_sq118 = xn3 & multm_reduce_sa128;
  assign multm_reduce_mulsc_mulb_sq119 = xn3 & multm_reduce_sa129;
  assign multm_reduce_mulsc_mulb_sq120 = xn3 & multm_reduce_sa130;
  assign multm_reduce_mulsc_mulb_sq121 = xn3 & multm_reduce_sa131;
  assign multm_reduce_mulsc_mulb_sq122 = xn3 & multm_reduce_sa132;
  assign multm_reduce_mulsc_mulb_sq123 = xn3 & multm_reduce_sa133;
  assign multm_reduce_mulsc_mulb_sq124 = xn3 & multm_reduce_sa134;
  assign multm_reduce_mulsc_mulb_sq125 = xn3 & multm_reduce_sa135;
  assign multm_reduce_mulsc_mulb_sq126 = xn3 & multm_reduce_sa136;
  assign multm_reduce_mulsc_mulb_sq127 = xn3 & multm_reduce_sa137;
  assign multm_reduce_mulsc_mulb_sq128 = xn3 & multm_reduce_sa138;
  assign multm_reduce_mulsc_mulb_sq129 = xn3 & multm_reduce_sa139;
  assign multm_reduce_mulsc_mulb_sq130 = xn3 & multm_reduce_sa140;
  assign multm_reduce_mulsc_mulb_sq131 = xn3 & multm_reduce_sa141;
  assign multm_reduce_mulsc_mulb_sq132 = xn3 & multm_reduce_sa142;
  assign multm_reduce_mulsc_mulb_sq133 = xn3 & multm_reduce_sa143;
  assign multm_reduce_mulsc_mulb_sq134 = xn3 & multm_reduce_sa144;
  assign multm_reduce_mulsc_mulb_sq135 = xn3 & multm_reduce_sa145;
  assign multm_reduce_mulsc_mulb_sq136 = xn3 & multm_reduce_sa146;
  assign multm_reduce_mulsc_mulb_sq137 = xn3 & multm_reduce_sa147;
  assign multm_reduce_mulsc_mulb_sq138 = xn3 & multm_reduce_sa148;
  assign multm_reduce_mulsc_mulb_sq139 = xn3 & multm_reduce_sa149;
  assign multm_reduce_mulsc_mulb_sq140 = xn3 & multm_reduce_sa150;
  assign multm_reduce_mulsc_mulb_sq141 = xn3 & multm_reduce_sa151;
  assign multm_reduce_mulsc_mulb_sq142 = xn3 & multm_reduce_sa152;
  assign multm_reduce_mulsc_mulb_sq143 = xn3 & multm_reduce_sa153;
  assign multm_reduce_mulsc_mulb_sq144 = xn3 & multm_reduce_sa154;
  assign multm_reduce_mulsc_mulb_sq145 = xn3 & multm_reduce_sa155;
  assign multm_reduce_mulsc_mulb_sq146 = xn3 & multm_reduce_sa156;
  assign multm_reduce_mulsc_mulb_sq147 = xn3 & multm_reduce_sa157;
  assign multm_reduce_mulsc_mulb_sq148 = xn3 & multm_reduce_sa158;
  assign multm_reduce_mulsc_mulb_sq149 = xn3 & multm_reduce_sa159;
  assign multm_reduce_mulsc_mulb_sq150 = xn3 & multm_reduce_sa160;
  assign multm_reduce_mulsc_mulb_sq151 = xn3 & multm_reduce_sa161;
  assign multm_reduce_mulsc_mulb_sq152 = xn3 & multm_reduce_sa162;
  assign multm_reduce_mulsc_mulb_sq153 = xn3 & multm_reduce_sa163;
  assign multm_reduce_mulsc_mulb_sq154 = xn3 & multm_reduce_sa164;
  assign multm_reduce_mulsc_mulb_sq155 = xn3 & multm_reduce_sa165;
  assign multm_reduce_mulsc_mulb_sq156 = xn3 & multm_reduce_sa166;
  assign multm_reduce_mulsc_mulb_sq157 = xn3 & multm_reduce_sa167;
  assign multm_reduce_mulsc_mulb_sq158 = xn3 & multm_reduce_sa168;
  assign multm_reduce_mulsc_mulb_sq159 = xn3 & multm_reduce_sa169;
  assign multm_reduce_mulsc_mulb_sq160 = xn3 & multm_reduce_sa170;
  assign multm_reduce_mulsc_mulb_sq161 = xn3 & multm_reduce_sa171;
  assign multm_reduce_mulsc_mulb_sq162 = xn3 & multm_reduce_sa172;
  assign multm_reduce_mulsc_mulb_sq163 = xn3 & multm_reduce_sa173;
  assign multm_reduce_mulsc_mulb_sq164 = xn3 & multm_reduce_sa174;
  assign multm_reduce_mulsc_mulb_sq165 = xn3 & multm_reduce_sa175;
  assign multm_reduce_mulsc_mulb_sq166 = xn3 & multm_reduce_sa176;
  assign multm_reduce_mulsc_mulb_sq167 = xn3 & multm_reduce_sa177;
  assign multm_reduce_mulsc_mulb_sq168 = xn3 & multm_reduce_sa178;
  assign multm_reduce_mulsc_mulb_sq169 = xn3 & multm_reduce_sa179;
  assign multm_reduce_mulsc_mulb_sq170 = xn3 & multm_reduce_sa180;
  assign multm_reduce_mulsc_mulb_sq171 = xn3 & multm_reduce_sa181;
  assign multm_reduce_mulsc_mulb_sq172 = xn3 & multm_reduce_sa182;
  assign multm_reduce_mulsc_mulb_sq173 = xn3 & multm_reduce_sa183;
  assign multm_reduce_mulsc_mulb_sq174 = xn3 & multm_reduce_sa184;
  assign multm_reduce_mulsc_mulb_sq175 = xn3 & multm_reduce_sa185;
  assign multm_reduce_mulsc_mulb_sq176 = xn3 & multm_reduce_mulsc_mulb_sp176;
  assign multm_reduce_mulsc_mulb_sq177 = xn3 & multm_reduce_mulsc_mulb_sp177;
  assign multm_reduce_mulsc_mulb_sq178 = xn3 & multm_reduce_mulsc_mulb_sp178;
  assign multm_reduce_mulsc_mulb_sq179 = xn3 & multm_reduce_mulsc_mulb_sp179;
  assign multm_reduce_mulsc_mulb_sq180 = xn3 & multm_reduce_mulsc_mulb_sp180;
  assign multm_reduce_mulsc_mulb_sq181 = xn3 & multm_reduce_mulsc_mulb_sp181;
  assign multm_reduce_mulsc_mulb_sq182 = xn3 & multm_reduce_mulsc_mulb_sp182;
  assign multm_reduce_mulsc_mulb_sq183 = xn3 & multm_reduce_mulsc_mulb_sp183;
  assign multm_reduce_mulsc_mulb_yoc0 = multm_reduce_mulsc_xbd & yc0_o;
  assign multm_reduce_mulsc_mulb_yoc1 = multm_reduce_mulsc_xbd & yc1_o;
  assign multm_reduce_mulsc_mulb_yoc2 = multm_reduce_mulsc_xbd & yc2_o;
  assign multm_reduce_mulsc_mulb_yoc3 = multm_reduce_mulsc_xbd & yc3_o;
  assign multm_reduce_mulsc_mulb_yoc4 = multm_reduce_mulsc_xbd & yc4_o;
  assign multm_reduce_mulsc_mulb_yoc5 = multm_reduce_mulsc_xbd & yc5_o;
  assign multm_reduce_mulsc_mulb_yoc6 = multm_reduce_mulsc_xbd & yc6_o;
  assign multm_reduce_mulsc_mulb_yoc7 = multm_reduce_mulsc_xbd & yc7_o;
  assign multm_reduce_mulsc_mulb_yoc8 = multm_reduce_mulsc_xbd & yc8_o;
  assign multm_reduce_mulsc_mulb_yoc9 = multm_reduce_mulsc_xbd & yc9_o;
  assign multm_reduce_mulsc_mulb_yoc10 = multm_reduce_mulsc_xbd & yc10_o;
  assign multm_reduce_mulsc_mulb_yoc11 = multm_reduce_mulsc_xbd & yc11_o;
  assign multm_reduce_mulsc_mulb_yoc12 = multm_reduce_mulsc_xbd & yc12_o;
  assign multm_reduce_mulsc_mulb_yoc13 = multm_reduce_mulsc_xbd & yc13_o;
  assign multm_reduce_mulsc_mulb_yoc14 = multm_reduce_mulsc_xbd & yc14_o;
  assign multm_reduce_mulsc_mulb_yoc15 = multm_reduce_mulsc_xbd & yc15_o;
  assign multm_reduce_mulsc_mulb_yoc16 = multm_reduce_mulsc_xbd & yc16_o;
  assign multm_reduce_mulsc_mulb_yoc17 = multm_reduce_mulsc_xbd & yc17_o;
  assign multm_reduce_mulsc_mulb_yoc18 = multm_reduce_mulsc_xbd & yc18_o;
  assign multm_reduce_mulsc_mulb_yoc19 = multm_reduce_mulsc_xbd & yc19_o;
  assign multm_reduce_mulsc_mulb_yoc20 = multm_reduce_mulsc_xbd & yc20_o;
  assign multm_reduce_mulsc_mulb_yoc21 = multm_reduce_mulsc_xbd & yc21_o;
  assign multm_reduce_mulsc_mulb_yoc22 = multm_reduce_mulsc_xbd & yc22_o;
  assign multm_reduce_mulsc_mulb_yoc23 = multm_reduce_mulsc_xbd & yc23_o;
  assign multm_reduce_mulsc_mulb_yoc24 = multm_reduce_mulsc_xbd & yc24_o;
  assign multm_reduce_mulsc_mulb_yoc25 = multm_reduce_mulsc_xbd & yc25_o;
  assign multm_reduce_mulsc_mulb_yoc26 = multm_reduce_mulsc_xbd & yc26_o;
  assign multm_reduce_mulsc_mulb_yoc27 = multm_reduce_mulsc_xbd & yc27_o;
  assign multm_reduce_mulsc_mulb_yoc28 = multm_reduce_mulsc_xbd & yc28_o;
  assign multm_reduce_mulsc_mulb_yoc29 = multm_reduce_mulsc_xbd & yc29_o;
  assign multm_reduce_mulsc_mulb_yoc30 = multm_reduce_mulsc_xbd & yc30_o;
  assign multm_reduce_mulsc_mulb_yoc31 = multm_reduce_mulsc_xbd & yc31_o;
  assign multm_reduce_mulsc_mulb_yoc32 = multm_reduce_mulsc_xbd & yc32_o;
  assign multm_reduce_mulsc_mulb_yoc33 = multm_reduce_mulsc_xbd & yc33_o;
  assign multm_reduce_mulsc_mulb_yoc34 = multm_reduce_mulsc_xbd & yc34_o;
  assign multm_reduce_mulsc_mulb_yoc35 = multm_reduce_mulsc_xbd & yc35_o;
  assign multm_reduce_mulsc_mulb_yoc36 = multm_reduce_mulsc_xbd & yc36_o;
  assign multm_reduce_mulsc_mulb_yoc37 = multm_reduce_mulsc_xbd & yc37_o;
  assign multm_reduce_mulsc_mulb_yoc38 = multm_reduce_mulsc_xbd & yc38_o;
  assign multm_reduce_mulsc_mulb_yoc39 = multm_reduce_mulsc_xbd & yc39_o;
  assign multm_reduce_mulsc_mulb_yoc40 = multm_reduce_mulsc_xbd & yc40_o;
  assign multm_reduce_mulsc_mulb_yoc41 = multm_reduce_mulsc_xbd & yc41_o;
  assign multm_reduce_mulsc_mulb_yoc42 = multm_reduce_mulsc_xbd & yc42_o;
  assign multm_reduce_mulsc_mulb_yoc43 = multm_reduce_mulsc_xbd & yc43_o;
  assign multm_reduce_mulsc_mulb_yoc44 = multm_reduce_mulsc_xbd & yc44_o;
  assign multm_reduce_mulsc_mulb_yoc45 = multm_reduce_mulsc_xbd & yc45_o;
  assign multm_reduce_mulsc_mulb_yoc46 = multm_reduce_mulsc_xbd & yc46_o;
  assign multm_reduce_mulsc_mulb_yoc47 = multm_reduce_mulsc_xbd & yc47_o;
  assign multm_reduce_mulsc_mulb_yoc48 = multm_reduce_mulsc_xbd & yc48_o;
  assign multm_reduce_mulsc_mulb_yoc49 = multm_reduce_mulsc_xbd & yc49_o;
  assign multm_reduce_mulsc_mulb_yoc50 = multm_reduce_mulsc_xbd & yc50_o;
  assign multm_reduce_mulsc_mulb_yoc51 = multm_reduce_mulsc_xbd & yc51_o;
  assign multm_reduce_mulsc_mulb_yoc52 = multm_reduce_mulsc_xbd & yc52_o;
  assign multm_reduce_mulsc_mulb_yoc53 = multm_reduce_mulsc_xbd & yc53_o;
  assign multm_reduce_mulsc_mulb_yoc54 = multm_reduce_mulsc_xbd & yc54_o;
  assign multm_reduce_mulsc_mulb_yoc55 = multm_reduce_mulsc_xbd & yc55_o;
  assign multm_reduce_mulsc_mulb_yoc56 = multm_reduce_mulsc_xbd & yc56_o;
  assign multm_reduce_mulsc_mulb_yoc57 = multm_reduce_mulsc_xbd & yc57_o;
  assign multm_reduce_mulsc_mulb_yoc58 = multm_reduce_mulsc_xbd & yc58_o;
  assign multm_reduce_mulsc_mulb_yoc59 = multm_reduce_mulsc_xbd & yc59_o;
  assign multm_reduce_mulsc_mulb_yoc60 = multm_reduce_mulsc_xbd & yc60_o;
  assign multm_reduce_mulsc_mulb_yoc61 = multm_reduce_mulsc_xbd & yc61_o;
  assign multm_reduce_mulsc_mulb_yoc62 = multm_reduce_mulsc_xbd & yc62_o;
  assign multm_reduce_mulsc_mulb_yoc63 = multm_reduce_mulsc_xbd & yc63_o;
  assign multm_reduce_mulsc_mulb_yoc64 = multm_reduce_mulsc_xbd & yc64_o;
  assign multm_reduce_mulsc_mulb_yoc65 = multm_reduce_mulsc_xbd & yc65_o;
  assign multm_reduce_mulsc_mulb_yoc66 = multm_reduce_mulsc_xbd & yc66_o;
  assign multm_reduce_mulsc_mulb_yoc67 = multm_reduce_mulsc_xbd & yc67_o;
  assign multm_reduce_mulsc_mulb_yoc68 = multm_reduce_mulsc_xbd & yc68_o;
  assign multm_reduce_mulsc_mulb_yoc69 = multm_reduce_mulsc_xbd & yc69_o;
  assign multm_reduce_mulsc_mulb_yoc70 = multm_reduce_mulsc_xbd & yc70_o;
  assign multm_reduce_mulsc_mulb_yoc71 = multm_reduce_mulsc_xbd & yc71_o;
  assign multm_reduce_mulsc_mulb_yoc72 = multm_reduce_mulsc_xbd & yc72_o;
  assign multm_reduce_mulsc_mulb_yoc73 = multm_reduce_mulsc_xbd & yc73_o;
  assign multm_reduce_mulsc_mulb_yoc74 = multm_reduce_mulsc_xbd & yc74_o;
  assign multm_reduce_mulsc_mulb_yoc75 = multm_reduce_mulsc_xbd & yc75_o;
  assign multm_reduce_mulsc_mulb_yoc76 = multm_reduce_mulsc_xbd & yc76_o;
  assign multm_reduce_mulsc_mulb_yoc77 = multm_reduce_mulsc_xbd & yc77_o;
  assign multm_reduce_mulsc_mulb_yoc78 = multm_reduce_mulsc_xbd & yc78_o;
  assign multm_reduce_mulsc_mulb_yoc79 = multm_reduce_mulsc_xbd & yc79_o;
  assign multm_reduce_mulsc_mulb_yoc80 = multm_reduce_mulsc_xbd & yc80_o;
  assign multm_reduce_mulsc_mulb_yoc81 = multm_reduce_mulsc_xbd & yc81_o;
  assign multm_reduce_mulsc_mulb_yoc82 = multm_reduce_mulsc_xbd & yc82_o;
  assign multm_reduce_mulsc_mulb_yoc83 = multm_reduce_mulsc_xbd & yc83_o;
  assign multm_reduce_mulsc_mulb_yoc84 = multm_reduce_mulsc_xbd & yc84_o;
  assign multm_reduce_mulsc_mulb_yoc85 = multm_reduce_mulsc_xbd & yc85_o;
  assign multm_reduce_mulsc_mulb_yoc86 = multm_reduce_mulsc_xbd & yc86_o;
  assign multm_reduce_mulsc_mulb_yoc87 = multm_reduce_mulsc_xbd & yc87_o;
  assign multm_reduce_mulsc_mulb_yoc88 = multm_reduce_mulsc_xbd & yc88_o;
  assign multm_reduce_mulsc_mulb_yoc89 = multm_reduce_mulsc_xbd & yc89_o;
  assign multm_reduce_mulsc_mulb_yoc90 = multm_reduce_mulsc_xbd & yc90_o;
  assign multm_reduce_mulsc_mulb_yoc91 = multm_reduce_mulsc_xbd & yc91_o;
  assign multm_reduce_mulsc_mulb_yoc92 = multm_reduce_mulsc_xbd & yc92_o;
  assign multm_reduce_mulsc_mulb_yoc93 = multm_reduce_mulsc_xbd & yc93_o;
  assign multm_reduce_mulsc_mulb_yoc94 = multm_reduce_mulsc_xbd & yc94_o;
  assign multm_reduce_mulsc_mulb_yoc95 = multm_reduce_mulsc_xbd & yc95_o;
  assign multm_reduce_mulsc_mulb_yoc96 = multm_reduce_mulsc_xbd & yc96_o;
  assign multm_reduce_mulsc_mulb_yoc97 = multm_reduce_mulsc_xbd & yc97_o;
  assign multm_reduce_mulsc_mulb_yoc98 = multm_reduce_mulsc_xbd & yc98_o;
  assign multm_reduce_mulsc_mulb_yoc99 = multm_reduce_mulsc_xbd & yc99_o;
  assign multm_reduce_mulsc_mulb_yoc100 = multm_reduce_mulsc_xbd & yc100_o;
  assign multm_reduce_mulsc_mulb_yoc101 = multm_reduce_mulsc_xbd & yc101_o;
  assign multm_reduce_mulsc_mulb_yoc102 = multm_reduce_mulsc_xbd & yc102_o;
  assign multm_reduce_mulsc_mulb_yoc103 = multm_reduce_mulsc_xbd & yc103_o;
  assign multm_reduce_mulsc_mulb_yoc104 = multm_reduce_mulsc_xbd & yc104_o;
  assign multm_reduce_mulsc_mulb_yoc105 = multm_reduce_mulsc_xbd & yc105_o;
  assign multm_reduce_mulsc_mulb_yoc106 = multm_reduce_mulsc_xbd & yc106_o;
  assign multm_reduce_mulsc_mulb_yoc107 = multm_reduce_mulsc_xbd & yc107_o;
  assign multm_reduce_mulsc_mulb_yoc108 = multm_reduce_mulsc_xbd & yc108_o;
  assign multm_reduce_mulsc_mulb_yoc109 = multm_reduce_mulsc_xbd & yc109_o;
  assign multm_reduce_mulsc_mulb_yoc110 = multm_reduce_mulsc_xbd & yc110_o;
  assign multm_reduce_mulsc_mulb_yoc111 = multm_reduce_mulsc_xbd & yc111_o;
  assign multm_reduce_mulsc_mulb_yoc112 = multm_reduce_mulsc_xbd & yc112_o;
  assign multm_reduce_mulsc_mulb_yoc113 = multm_reduce_mulsc_xbd & yc113_o;
  assign multm_reduce_mulsc_mulb_yoc114 = multm_reduce_mulsc_xbd & yc114_o;
  assign multm_reduce_mulsc_mulb_yoc115 = multm_reduce_mulsc_xbd & yc115_o;
  assign multm_reduce_mulsc_mulb_yoc116 = multm_reduce_mulsc_xbd & yc116_o;
  assign multm_reduce_mulsc_mulb_yoc117 = multm_reduce_mulsc_xbd & yc117_o;
  assign multm_reduce_mulsc_mulb_yoc118 = multm_reduce_mulsc_xbd & yc118_o;
  assign multm_reduce_mulsc_mulb_yoc119 = multm_reduce_mulsc_xbd & yc119_o;
  assign multm_reduce_mulsc_mulb_yoc120 = multm_reduce_mulsc_xbd & yc120_o;
  assign multm_reduce_mulsc_mulb_yoc121 = multm_reduce_mulsc_xbd & yc121_o;
  assign multm_reduce_mulsc_mulb_yoc122 = multm_reduce_mulsc_xbd & yc122_o;
  assign multm_reduce_mulsc_mulb_yoc123 = multm_reduce_mulsc_xbd & yc123_o;
  assign multm_reduce_mulsc_mulb_yoc124 = multm_reduce_mulsc_xbd & yc124_o;
  assign multm_reduce_mulsc_mulb_yoc125 = multm_reduce_mulsc_xbd & yc125_o;
  assign multm_reduce_mulsc_mulb_yoc126 = multm_reduce_mulsc_xbd & yc126_o;
  assign multm_reduce_mulsc_mulb_yoc127 = multm_reduce_mulsc_xbd & yc127_o;
  assign multm_reduce_mulsc_mulb_yoc128 = multm_reduce_mulsc_xbd & yc128_o;
  assign multm_reduce_mulsc_mulb_yoc129 = multm_reduce_mulsc_xbd & yc129_o;
  assign multm_reduce_mulsc_mulb_yoc130 = multm_reduce_mulsc_xbd & yc130_o;
  assign multm_reduce_mulsc_mulb_yoc131 = multm_reduce_mulsc_xbd & yc131_o;
  assign multm_reduce_mulsc_mulb_yoc132 = multm_reduce_mulsc_xbd & yc132_o;
  assign multm_reduce_mulsc_mulb_yoc133 = multm_reduce_mulsc_xbd & yc133_o;
  assign multm_reduce_mulsc_mulb_yoc134 = multm_reduce_mulsc_xbd & yc134_o;
  assign multm_reduce_mulsc_mulb_yoc135 = multm_reduce_mulsc_xbd & yc135_o;
  assign multm_reduce_mulsc_mulb_yoc136 = multm_reduce_mulsc_xbd & yc136_o;
  assign multm_reduce_mulsc_mulb_yoc137 = multm_reduce_mulsc_xbd & yc137_o;
  assign multm_reduce_mulsc_mulb_yoc138 = multm_reduce_mulsc_xbd & yc138_o;
  assign multm_reduce_mulsc_mulb_yoc139 = multm_reduce_mulsc_xbd & yc139_o;
  assign multm_reduce_mulsc_mulb_yoc140 = multm_reduce_mulsc_xbd & yc140_o;
  assign multm_reduce_mulsc_mulb_yoc141 = multm_reduce_mulsc_xbd & yc141_o;
  assign multm_reduce_mulsc_mulb_yoc142 = multm_reduce_mulsc_xbd & yc142_o;
  assign multm_reduce_mulsc_mulb_yoc143 = multm_reduce_mulsc_xbd & yc143_o;
  assign multm_reduce_mulsc_mulb_yoc144 = multm_reduce_mulsc_xbd & yc144_o;
  assign multm_reduce_mulsc_mulb_yoc145 = multm_reduce_mulsc_xbd & yc145_o;
  assign multm_reduce_mulsc_mulb_yoc146 = multm_reduce_mulsc_xbd & yc146_o;
  assign multm_reduce_mulsc_mulb_yoc147 = multm_reduce_mulsc_xbd & yc147_o;
  assign multm_reduce_mulsc_mulb_yoc148 = multm_reduce_mulsc_xbd & yc148_o;
  assign multm_reduce_mulsc_mulb_yoc149 = multm_reduce_mulsc_xbd & yc149_o;
  assign multm_reduce_mulsc_mulb_yoc150 = multm_reduce_mulsc_xbd & yc150_o;
  assign multm_reduce_mulsc_mulb_yoc151 = multm_reduce_mulsc_xbd & yc151_o;
  assign multm_reduce_mulsc_mulb_yoc152 = multm_reduce_mulsc_xbd & yc152_o;
  assign multm_reduce_mulsc_mulb_yoc153 = multm_reduce_mulsc_xbd & yc153_o;
  assign multm_reduce_mulsc_mulb_yoc154 = multm_reduce_mulsc_xbd & yc154_o;
  assign multm_reduce_mulsc_mulb_yoc155 = multm_reduce_mulsc_xbd & yc155_o;
  assign multm_reduce_mulsc_mulb_yoc156 = multm_reduce_mulsc_xbd & yc156_o;
  assign multm_reduce_mulsc_mulb_yoc157 = multm_reduce_mulsc_xbd & yc157_o;
  assign multm_reduce_mulsc_mulb_yoc158 = multm_reduce_mulsc_xbd & yc158_o;
  assign multm_reduce_mulsc_mulb_yoc159 = multm_reduce_mulsc_xbd & yc159_o;
  assign multm_reduce_mulsc_mulb_yoc160 = multm_reduce_mulsc_xbd & yc160_o;
  assign multm_reduce_mulsc_mulb_yoc161 = multm_reduce_mulsc_xbd & yc161_o;
  assign multm_reduce_mulsc_mulb_yoc162 = multm_reduce_mulsc_xbd & yc162_o;
  assign multm_reduce_mulsc_mulb_yoc163 = multm_reduce_mulsc_xbd & yc163_o;
  assign multm_reduce_mulsc_mulb_yoc164 = multm_reduce_mulsc_xbd & yc164_o;
  assign multm_reduce_mulsc_mulb_yoc165 = multm_reduce_mulsc_xbd & yc165_o;
  assign multm_reduce_mulsc_mulb_yoc166 = multm_reduce_mulsc_xbd & yc166_o;
  assign multm_reduce_mulsc_mulb_yoc167 = multm_reduce_mulsc_xbd & yc167_o;
  assign multm_reduce_mulsc_mulb_yoc168 = multm_reduce_mulsc_xbd & yc168_o;
  assign multm_reduce_mulsc_mulb_yoc169 = multm_reduce_mulsc_xbd & yc169_o;
  assign multm_reduce_mulsc_mulb_yoc170 = multm_reduce_mulsc_xbd & yc170_o;
  assign multm_reduce_mulsc_mulb_yoc171 = multm_reduce_mulsc_xbd & yc171_o;
  assign multm_reduce_mulsc_mulb_yoc172 = multm_reduce_mulsc_xbd & yc172_o;
  assign multm_reduce_mulsc_mulb_yoc173 = multm_reduce_mulsc_xbd & yc173_o;
  assign multm_reduce_mulsc_mulb_yoc174 = multm_reduce_mulsc_xbd & yc174_o;
  assign multm_reduce_mulsc_mulb_yoc175 = multm_reduce_mulsc_xbd & yc175_o;
  assign multm_reduce_mulsc_mulb_yoc176 = multm_reduce_mulsc_xbd & yc176_o;
  assign multm_reduce_mulsc_mulb_yoc177 = multm_reduce_mulsc_xbd & yc177_o;
  assign multm_reduce_mulsc_mulb_yoc178 = multm_reduce_mulsc_xbd & yc178_o;
  assign multm_reduce_mulsc_mulb_yoc179 = multm_reduce_mulsc_xbd & yc179_o;
  assign multm_reduce_mulsc_mulb_yoc180 = multm_reduce_mulsc_xbd & yc180_o;
  assign multm_reduce_mulsc_mulb_yoc181 = multm_reduce_mulsc_xbd & yc181_o;
  assign multm_reduce_mulsc_mulb_yoc182 = multm_reduce_mulsc_xbd & yc182_o;
  assign multm_reduce_mulsc_mulb_yoc183 = multm_reduce_mulsc_xbd & yc183_o;
  assign multm_reduce_mulsc_mulb_yos0 = multm_reduce_mulsc_xbd & ys0_o;
  assign multm_reduce_mulsc_mulb_yos1 = multm_reduce_mulsc_xbd & ys1_o;
  assign multm_reduce_mulsc_mulb_yos2 = multm_reduce_mulsc_xbd & ys2_o;
  assign multm_reduce_mulsc_mulb_yos3 = multm_reduce_mulsc_xbd & ys3_o;
  assign multm_reduce_mulsc_mulb_yos4 = multm_reduce_mulsc_xbd & ys4_o;
  assign multm_reduce_mulsc_mulb_yos5 = multm_reduce_mulsc_xbd & ys5_o;
  assign multm_reduce_mulsc_mulb_yos6 = multm_reduce_mulsc_xbd & ys6_o;
  assign multm_reduce_mulsc_mulb_yos7 = multm_reduce_mulsc_xbd & ys7_o;
  assign multm_reduce_mulsc_mulb_yos8 = multm_reduce_mulsc_xbd & ys8_o;
  assign multm_reduce_mulsc_mulb_yos9 = multm_reduce_mulsc_xbd & ys9_o;
  assign multm_reduce_mulsc_mulb_yos10 = multm_reduce_mulsc_xbd & ys10_o;
  assign multm_reduce_mulsc_mulb_yos11 = multm_reduce_mulsc_xbd & ys11_o;
  assign multm_reduce_mulsc_mulb_yos12 = multm_reduce_mulsc_xbd & ys12_o;
  assign multm_reduce_mulsc_mulb_yos13 = multm_reduce_mulsc_xbd & ys13_o;
  assign multm_reduce_mulsc_mulb_yos14 = multm_reduce_mulsc_xbd & ys14_o;
  assign multm_reduce_mulsc_mulb_yos15 = multm_reduce_mulsc_xbd & ys15_o;
  assign multm_reduce_mulsc_mulb_yos16 = multm_reduce_mulsc_xbd & ys16_o;
  assign multm_reduce_mulsc_mulb_yos17 = multm_reduce_mulsc_xbd & ys17_o;
  assign multm_reduce_mulsc_mulb_yos18 = multm_reduce_mulsc_xbd & ys18_o;
  assign multm_reduce_mulsc_mulb_yos19 = multm_reduce_mulsc_xbd & ys19_o;
  assign multm_reduce_mulsc_mulb_yos20 = multm_reduce_mulsc_xbd & ys20_o;
  assign multm_reduce_mulsc_mulb_yos21 = multm_reduce_mulsc_xbd & ys21_o;
  assign multm_reduce_mulsc_mulb_yos22 = multm_reduce_mulsc_xbd & ys22_o;
  assign multm_reduce_mulsc_mulb_yos23 = multm_reduce_mulsc_xbd & ys23_o;
  assign multm_reduce_mulsc_mulb_yos24 = multm_reduce_mulsc_xbd & ys24_o;
  assign multm_reduce_mulsc_mulb_yos25 = multm_reduce_mulsc_xbd & ys25_o;
  assign multm_reduce_mulsc_mulb_yos26 = multm_reduce_mulsc_xbd & ys26_o;
  assign multm_reduce_mulsc_mulb_yos27 = multm_reduce_mulsc_xbd & ys27_o;
  assign multm_reduce_mulsc_mulb_yos28 = multm_reduce_mulsc_xbd & ys28_o;
  assign multm_reduce_mulsc_mulb_yos29 = multm_reduce_mulsc_xbd & ys29_o;
  assign multm_reduce_mulsc_mulb_yos30 = multm_reduce_mulsc_xbd & ys30_o;
  assign multm_reduce_mulsc_mulb_yos31 = multm_reduce_mulsc_xbd & ys31_o;
  assign multm_reduce_mulsc_mulb_yos32 = multm_reduce_mulsc_xbd & ys32_o;
  assign multm_reduce_mulsc_mulb_yos33 = multm_reduce_mulsc_xbd & ys33_o;
  assign multm_reduce_mulsc_mulb_yos34 = multm_reduce_mulsc_xbd & ys34_o;
  assign multm_reduce_mulsc_mulb_yos35 = multm_reduce_mulsc_xbd & ys35_o;
  assign multm_reduce_mulsc_mulb_yos36 = multm_reduce_mulsc_xbd & ys36_o;
  assign multm_reduce_mulsc_mulb_yos37 = multm_reduce_mulsc_xbd & ys37_o;
  assign multm_reduce_mulsc_mulb_yos38 = multm_reduce_mulsc_xbd & ys38_o;
  assign multm_reduce_mulsc_mulb_yos39 = multm_reduce_mulsc_xbd & ys39_o;
  assign multm_reduce_mulsc_mulb_yos40 = multm_reduce_mulsc_xbd & ys40_o;
  assign multm_reduce_mulsc_mulb_yos41 = multm_reduce_mulsc_xbd & ys41_o;
  assign multm_reduce_mulsc_mulb_yos42 = multm_reduce_mulsc_xbd & ys42_o;
  assign multm_reduce_mulsc_mulb_yos43 = multm_reduce_mulsc_xbd & ys43_o;
  assign multm_reduce_mulsc_mulb_yos44 = multm_reduce_mulsc_xbd & ys44_o;
  assign multm_reduce_mulsc_mulb_yos45 = multm_reduce_mulsc_xbd & ys45_o;
  assign multm_reduce_mulsc_mulb_yos46 = multm_reduce_mulsc_xbd & ys46_o;
  assign multm_reduce_mulsc_mulb_yos47 = multm_reduce_mulsc_xbd & ys47_o;
  assign multm_reduce_mulsc_mulb_yos48 = multm_reduce_mulsc_xbd & ys48_o;
  assign multm_reduce_mulsc_mulb_yos49 = multm_reduce_mulsc_xbd & ys49_o;
  assign multm_reduce_mulsc_mulb_yos50 = multm_reduce_mulsc_xbd & ys50_o;
  assign multm_reduce_mulsc_mulb_yos51 = multm_reduce_mulsc_xbd & ys51_o;
  assign multm_reduce_mulsc_mulb_yos52 = multm_reduce_mulsc_xbd & ys52_o;
  assign multm_reduce_mulsc_mulb_yos53 = multm_reduce_mulsc_xbd & ys53_o;
  assign multm_reduce_mulsc_mulb_yos54 = multm_reduce_mulsc_xbd & ys54_o;
  assign multm_reduce_mulsc_mulb_yos55 = multm_reduce_mulsc_xbd & ys55_o;
  assign multm_reduce_mulsc_mulb_yos56 = multm_reduce_mulsc_xbd & ys56_o;
  assign multm_reduce_mulsc_mulb_yos57 = multm_reduce_mulsc_xbd & ys57_o;
  assign multm_reduce_mulsc_mulb_yos58 = multm_reduce_mulsc_xbd & ys58_o;
  assign multm_reduce_mulsc_mulb_yos59 = multm_reduce_mulsc_xbd & ys59_o;
  assign multm_reduce_mulsc_mulb_yos60 = multm_reduce_mulsc_xbd & ys60_o;
  assign multm_reduce_mulsc_mulb_yos61 = multm_reduce_mulsc_xbd & ys61_o;
  assign multm_reduce_mulsc_mulb_yos62 = multm_reduce_mulsc_xbd & ys62_o;
  assign multm_reduce_mulsc_mulb_yos63 = multm_reduce_mulsc_xbd & ys63_o;
  assign multm_reduce_mulsc_mulb_yos64 = multm_reduce_mulsc_xbd & ys64_o;
  assign multm_reduce_mulsc_mulb_yos65 = multm_reduce_mulsc_xbd & ys65_o;
  assign multm_reduce_mulsc_mulb_yos66 = multm_reduce_mulsc_xbd & ys66_o;
  assign multm_reduce_mulsc_mulb_yos67 = multm_reduce_mulsc_xbd & ys67_o;
  assign multm_reduce_mulsc_mulb_yos68 = multm_reduce_mulsc_xbd & ys68_o;
  assign multm_reduce_mulsc_mulb_yos69 = multm_reduce_mulsc_xbd & ys69_o;
  assign multm_reduce_mulsc_mulb_yos70 = multm_reduce_mulsc_xbd & ys70_o;
  assign multm_reduce_mulsc_mulb_yos71 = multm_reduce_mulsc_xbd & ys71_o;
  assign multm_reduce_mulsc_mulb_yos72 = multm_reduce_mulsc_xbd & ys72_o;
  assign multm_reduce_mulsc_mulb_yos73 = multm_reduce_mulsc_xbd & ys73_o;
  assign multm_reduce_mulsc_mulb_yos74 = multm_reduce_mulsc_xbd & ys74_o;
  assign multm_reduce_mulsc_mulb_yos75 = multm_reduce_mulsc_xbd & ys75_o;
  assign multm_reduce_mulsc_mulb_yos76 = multm_reduce_mulsc_xbd & ys76_o;
  assign multm_reduce_mulsc_mulb_yos77 = multm_reduce_mulsc_xbd & ys77_o;
  assign multm_reduce_mulsc_mulb_yos78 = multm_reduce_mulsc_xbd & ys78_o;
  assign multm_reduce_mulsc_mulb_yos79 = multm_reduce_mulsc_xbd & ys79_o;
  assign multm_reduce_mulsc_mulb_yos80 = multm_reduce_mulsc_xbd & ys80_o;
  assign multm_reduce_mulsc_mulb_yos81 = multm_reduce_mulsc_xbd & ys81_o;
  assign multm_reduce_mulsc_mulb_yos82 = multm_reduce_mulsc_xbd & ys82_o;
  assign multm_reduce_mulsc_mulb_yos83 = multm_reduce_mulsc_xbd & ys83_o;
  assign multm_reduce_mulsc_mulb_yos84 = multm_reduce_mulsc_xbd & ys84_o;
  assign multm_reduce_mulsc_mulb_yos85 = multm_reduce_mulsc_xbd & ys85_o;
  assign multm_reduce_mulsc_mulb_yos86 = multm_reduce_mulsc_xbd & ys86_o;
  assign multm_reduce_mulsc_mulb_yos87 = multm_reduce_mulsc_xbd & ys87_o;
  assign multm_reduce_mulsc_mulb_yos88 = multm_reduce_mulsc_xbd & ys88_o;
  assign multm_reduce_mulsc_mulb_yos89 = multm_reduce_mulsc_xbd & ys89_o;
  assign multm_reduce_mulsc_mulb_yos90 = multm_reduce_mulsc_xbd & ys90_o;
  assign multm_reduce_mulsc_mulb_yos91 = multm_reduce_mulsc_xbd & ys91_o;
  assign multm_reduce_mulsc_mulb_yos92 = multm_reduce_mulsc_xbd & ys92_o;
  assign multm_reduce_mulsc_mulb_yos93 = multm_reduce_mulsc_xbd & ys93_o;
  assign multm_reduce_mulsc_mulb_yos94 = multm_reduce_mulsc_xbd & ys94_o;
  assign multm_reduce_mulsc_mulb_yos95 = multm_reduce_mulsc_xbd & ys95_o;
  assign multm_reduce_mulsc_mulb_yos96 = multm_reduce_mulsc_xbd & ys96_o;
  assign multm_reduce_mulsc_mulb_yos97 = multm_reduce_mulsc_xbd & ys97_o;
  assign multm_reduce_mulsc_mulb_yos98 = multm_reduce_mulsc_xbd & ys98_o;
  assign multm_reduce_mulsc_mulb_yos99 = multm_reduce_mulsc_xbd & ys99_o;
  assign multm_reduce_mulsc_mulb_yos100 = multm_reduce_mulsc_xbd & ys100_o;
  assign multm_reduce_mulsc_mulb_yos101 = multm_reduce_mulsc_xbd & ys101_o;
  assign multm_reduce_mulsc_mulb_yos102 = multm_reduce_mulsc_xbd & ys102_o;
  assign multm_reduce_mulsc_mulb_yos103 = multm_reduce_mulsc_xbd & ys103_o;
  assign multm_reduce_mulsc_mulb_yos104 = multm_reduce_mulsc_xbd & ys104_o;
  assign multm_reduce_mulsc_mulb_yos105 = multm_reduce_mulsc_xbd & ys105_o;
  assign multm_reduce_mulsc_mulb_yos106 = multm_reduce_mulsc_xbd & ys106_o;
  assign multm_reduce_mulsc_mulb_yos107 = multm_reduce_mulsc_xbd & ys107_o;
  assign multm_reduce_mulsc_mulb_yos108 = multm_reduce_mulsc_xbd & ys108_o;
  assign multm_reduce_mulsc_mulb_yos109 = multm_reduce_mulsc_xbd & ys109_o;
  assign multm_reduce_mulsc_mulb_yos110 = multm_reduce_mulsc_xbd & ys110_o;
  assign multm_reduce_mulsc_mulb_yos111 = multm_reduce_mulsc_xbd & ys111_o;
  assign multm_reduce_mulsc_mulb_yos112 = multm_reduce_mulsc_xbd & ys112_o;
  assign multm_reduce_mulsc_mulb_yos113 = multm_reduce_mulsc_xbd & ys113_o;
  assign multm_reduce_mulsc_mulb_yos114 = multm_reduce_mulsc_xbd & ys114_o;
  assign multm_reduce_mulsc_mulb_yos115 = multm_reduce_mulsc_xbd & ys115_o;
  assign multm_reduce_mulsc_mulb_yos116 = multm_reduce_mulsc_xbd & ys116_o;
  assign multm_reduce_mulsc_mulb_yos117 = multm_reduce_mulsc_xbd & ys117_o;
  assign multm_reduce_mulsc_mulb_yos118 = multm_reduce_mulsc_xbd & ys118_o;
  assign multm_reduce_mulsc_mulb_yos119 = multm_reduce_mulsc_xbd & ys119_o;
  assign multm_reduce_mulsc_mulb_yos120 = multm_reduce_mulsc_xbd & ys120_o;
  assign multm_reduce_mulsc_mulb_yos121 = multm_reduce_mulsc_xbd & ys121_o;
  assign multm_reduce_mulsc_mulb_yos122 = multm_reduce_mulsc_xbd & ys122_o;
  assign multm_reduce_mulsc_mulb_yos123 = multm_reduce_mulsc_xbd & ys123_o;
  assign multm_reduce_mulsc_mulb_yos124 = multm_reduce_mulsc_xbd & ys124_o;
  assign multm_reduce_mulsc_mulb_yos125 = multm_reduce_mulsc_xbd & ys125_o;
  assign multm_reduce_mulsc_mulb_yos126 = multm_reduce_mulsc_xbd & ys126_o;
  assign multm_reduce_mulsc_mulb_yos127 = multm_reduce_mulsc_xbd & ys127_o;
  assign multm_reduce_mulsc_mulb_yos128 = multm_reduce_mulsc_xbd & ys128_o;
  assign multm_reduce_mulsc_mulb_yos129 = multm_reduce_mulsc_xbd & ys129_o;
  assign multm_reduce_mulsc_mulb_yos130 = multm_reduce_mulsc_xbd & ys130_o;
  assign multm_reduce_mulsc_mulb_yos131 = multm_reduce_mulsc_xbd & ys131_o;
  assign multm_reduce_mulsc_mulb_yos132 = multm_reduce_mulsc_xbd & ys132_o;
  assign multm_reduce_mulsc_mulb_yos133 = multm_reduce_mulsc_xbd & ys133_o;
  assign multm_reduce_mulsc_mulb_yos134 = multm_reduce_mulsc_xbd & ys134_o;
  assign multm_reduce_mulsc_mulb_yos135 = multm_reduce_mulsc_xbd & ys135_o;
  assign multm_reduce_mulsc_mulb_yos136 = multm_reduce_mulsc_xbd & ys136_o;
  assign multm_reduce_mulsc_mulb_yos137 = multm_reduce_mulsc_xbd & ys137_o;
  assign multm_reduce_mulsc_mulb_yos138 = multm_reduce_mulsc_xbd & ys138_o;
  assign multm_reduce_mulsc_mulb_yos139 = multm_reduce_mulsc_xbd & ys139_o;
  assign multm_reduce_mulsc_mulb_yos140 = multm_reduce_mulsc_xbd & ys140_o;
  assign multm_reduce_mulsc_mulb_yos141 = multm_reduce_mulsc_xbd & ys141_o;
  assign multm_reduce_mulsc_mulb_yos142 = multm_reduce_mulsc_xbd & ys142_o;
  assign multm_reduce_mulsc_mulb_yos143 = multm_reduce_mulsc_xbd & ys143_o;
  assign multm_reduce_mulsc_mulb_yos144 = multm_reduce_mulsc_xbd & ys144_o;
  assign multm_reduce_mulsc_mulb_yos145 = multm_reduce_mulsc_xbd & ys145_o;
  assign multm_reduce_mulsc_mulb_yos146 = multm_reduce_mulsc_xbd & ys146_o;
  assign multm_reduce_mulsc_mulb_yos147 = multm_reduce_mulsc_xbd & ys147_o;
  assign multm_reduce_mulsc_mulb_yos148 = multm_reduce_mulsc_xbd & ys148_o;
  assign multm_reduce_mulsc_mulb_yos149 = multm_reduce_mulsc_xbd & ys149_o;
  assign multm_reduce_mulsc_mulb_yos150 = multm_reduce_mulsc_xbd & ys150_o;
  assign multm_reduce_mulsc_mulb_yos151 = multm_reduce_mulsc_xbd & ys151_o;
  assign multm_reduce_mulsc_mulb_yos152 = multm_reduce_mulsc_xbd & ys152_o;
  assign multm_reduce_mulsc_mulb_yos153 = multm_reduce_mulsc_xbd & ys153_o;
  assign multm_reduce_mulsc_mulb_yos154 = multm_reduce_mulsc_xbd & ys154_o;
  assign multm_reduce_mulsc_mulb_yos155 = multm_reduce_mulsc_xbd & ys155_o;
  assign multm_reduce_mulsc_mulb_yos156 = multm_reduce_mulsc_xbd & ys156_o;
  assign multm_reduce_mulsc_mulb_yos157 = multm_reduce_mulsc_xbd & ys157_o;
  assign multm_reduce_mulsc_mulb_yos158 = multm_reduce_mulsc_xbd & ys158_o;
  assign multm_reduce_mulsc_mulb_yos159 = multm_reduce_mulsc_xbd & ys159_o;
  assign multm_reduce_mulsc_mulb_yos160 = multm_reduce_mulsc_xbd & ys160_o;
  assign multm_reduce_mulsc_mulb_yos161 = multm_reduce_mulsc_xbd & ys161_o;
  assign multm_reduce_mulsc_mulb_yos162 = multm_reduce_mulsc_xbd & ys162_o;
  assign multm_reduce_mulsc_mulb_yos163 = multm_reduce_mulsc_xbd & ys163_o;
  assign multm_reduce_mulsc_mulb_yos164 = multm_reduce_mulsc_xbd & ys164_o;
  assign multm_reduce_mulsc_mulb_yos165 = multm_reduce_mulsc_xbd & ys165_o;
  assign multm_reduce_mulsc_mulb_yos166 = multm_reduce_mulsc_xbd & ys166_o;
  assign multm_reduce_mulsc_mulb_yos167 = multm_reduce_mulsc_xbd & ys167_o;
  assign multm_reduce_mulsc_mulb_yos168 = multm_reduce_mulsc_xbd & ys168_o;
  assign multm_reduce_mulsc_mulb_yos169 = multm_reduce_mulsc_xbd & ys169_o;
  assign multm_reduce_mulsc_mulb_yos170 = multm_reduce_mulsc_xbd & ys170_o;
  assign multm_reduce_mulsc_mulb_yos171 = multm_reduce_mulsc_xbd & ys171_o;
  assign multm_reduce_mulsc_mulb_yos172 = multm_reduce_mulsc_xbd & ys172_o;
  assign multm_reduce_mulsc_mulb_yos173 = multm_reduce_mulsc_xbd & ys173_o;
  assign multm_reduce_mulsc_mulb_yos174 = multm_reduce_mulsc_xbd & ys174_o;
  assign multm_reduce_mulsc_mulb_yos175 = multm_reduce_mulsc_xbd & ys175_o;
  assign multm_reduce_mulsc_mulb_yos176 = multm_reduce_mulsc_xbd & ys176_o;
  assign multm_reduce_mulsc_mulb_yos177 = multm_reduce_mulsc_xbd & ys177_o;
  assign multm_reduce_mulsc_mulb_yos178 = multm_reduce_mulsc_xbd & ys178_o;
  assign multm_reduce_mulsc_mulb_yos179 = multm_reduce_mulsc_xbd & ys179_o;
  assign multm_reduce_mulsc_mulb_yos180 = multm_reduce_mulsc_xbd & ys180_o;
  assign multm_reduce_mulsc_mulb_yos181 = multm_reduce_mulsc_xbd & ys181_o;
  assign multm_reduce_mulsc_mulb_yos182 = multm_reduce_mulsc_xbd & ys182_o;
  assign multm_reduce_mulsc_mulb_yos183 = multm_reduce_mulsc_xbd & ys183_o;
  assign multm_reduce_mulsc_shrsc_cq0 = multm_reduce_mulsc_shrsc_sp0 & multm_reduce_mulsc_shrsc_cp0;
  assign multm_reduce_mulsc_shrsc_cq1 = multm_reduce_mulsc_shrsc_sp1 & multm_reduce_mulsc_shrsc_cp1;
  assign multm_reduce_mulsc_shrsc_cq2 = multm_reduce_mulsc_shrsc_sp2 & multm_reduce_mulsc_shrsc_cp2;
  assign multm_reduce_mulsc_shrsc_cq3 = multm_reduce_mulsc_shrsc_sp3 & multm_reduce_mulsc_shrsc_cp3;
  assign multm_reduce_mulsc_shrsc_cq4 = multm_reduce_mulsc_shrsc_sp4 & multm_reduce_mulsc_shrsc_cp4;
  assign multm_reduce_mulsc_shrsc_cq5 = multm_reduce_mulsc_shrsc_sp5 & multm_reduce_mulsc_shrsc_cp5;
  assign multm_reduce_mulsc_shrsc_cq6 = multm_reduce_mulsc_shrsc_sp6 & multm_reduce_mulsc_shrsc_cp6;
  assign multm_reduce_mulsc_shrsc_cq7 = multm_reduce_mulsc_shrsc_sp7 & multm_reduce_mulsc_shrsc_cp7;
  assign multm_reduce_mulsc_shrsc_cq8 = multm_reduce_mulsc_shrsc_sp8 & multm_reduce_mulsc_shrsc_cp8;
  assign multm_reduce_mulsc_shrsc_cq9 = multm_reduce_mulsc_shrsc_sp9 & multm_reduce_mulsc_shrsc_cp9;
  assign multm_reduce_mulsc_shrsc_cq10 = multm_reduce_mulsc_shrsc_sp10 & multm_reduce_mulsc_shrsc_cp10;
  assign multm_reduce_mulsc_shrsc_cq11 = multm_reduce_mulsc_shrsc_sp11 & multm_reduce_mulsc_shrsc_cp11;
  assign multm_reduce_mulsc_shrsc_cq12 = multm_reduce_mulsc_shrsc_sp12 & multm_reduce_mulsc_shrsc_cp12;
  assign multm_reduce_mulsc_shrsc_cq13 = multm_reduce_mulsc_shrsc_sp13 & multm_reduce_mulsc_shrsc_cp13;
  assign multm_reduce_mulsc_shrsc_cq14 = multm_reduce_mulsc_shrsc_sp14 & multm_reduce_mulsc_shrsc_cp14;
  assign multm_reduce_mulsc_shrsc_cq15 = multm_reduce_mulsc_shrsc_sp15 & multm_reduce_mulsc_shrsc_cp15;
  assign multm_reduce_mulsc_shrsc_cq16 = multm_reduce_mulsc_shrsc_sp16 & multm_reduce_mulsc_shrsc_cp16;
  assign multm_reduce_mulsc_shrsc_cq17 = multm_reduce_mulsc_shrsc_sp17 & multm_reduce_mulsc_shrsc_cp17;
  assign multm_reduce_mulsc_shrsc_cq18 = multm_reduce_mulsc_shrsc_sp18 & multm_reduce_mulsc_shrsc_cp18;
  assign multm_reduce_mulsc_shrsc_cq19 = multm_reduce_mulsc_shrsc_sp19 & multm_reduce_mulsc_shrsc_cp19;
  assign multm_reduce_mulsc_shrsc_cq20 = multm_reduce_mulsc_shrsc_sp20 & multm_reduce_mulsc_shrsc_cp20;
  assign multm_reduce_mulsc_shrsc_cq21 = multm_reduce_mulsc_shrsc_sp21 & multm_reduce_mulsc_shrsc_cp21;
  assign multm_reduce_mulsc_shrsc_cq22 = multm_reduce_mulsc_shrsc_sp22 & multm_reduce_mulsc_shrsc_cp22;
  assign multm_reduce_mulsc_shrsc_cq23 = multm_reduce_mulsc_shrsc_sp23 & multm_reduce_mulsc_shrsc_cp23;
  assign multm_reduce_mulsc_shrsc_cq24 = multm_reduce_mulsc_shrsc_sp24 & multm_reduce_mulsc_shrsc_cp24;
  assign multm_reduce_mulsc_shrsc_cq25 = multm_reduce_mulsc_shrsc_sp25 & multm_reduce_mulsc_shrsc_cp25;
  assign multm_reduce_mulsc_shrsc_cq26 = multm_reduce_mulsc_shrsc_sp26 & multm_reduce_mulsc_shrsc_cp26;
  assign multm_reduce_mulsc_shrsc_cq27 = multm_reduce_mulsc_shrsc_sp27 & multm_reduce_mulsc_shrsc_cp27;
  assign multm_reduce_mulsc_shrsc_cq28 = multm_reduce_mulsc_shrsc_sp28 & multm_reduce_mulsc_shrsc_cp28;
  assign multm_reduce_mulsc_shrsc_cq29 = multm_reduce_mulsc_shrsc_sp29 & multm_reduce_mulsc_shrsc_cp29;
  assign multm_reduce_mulsc_shrsc_cq30 = multm_reduce_mulsc_shrsc_sp30 & multm_reduce_mulsc_shrsc_cp30;
  assign multm_reduce_mulsc_shrsc_cq31 = multm_reduce_mulsc_shrsc_sp31 & multm_reduce_mulsc_shrsc_cp31;
  assign multm_reduce_mulsc_shrsc_cq32 = multm_reduce_mulsc_shrsc_sp32 & multm_reduce_mulsc_shrsc_cp32;
  assign multm_reduce_mulsc_shrsc_cq33 = multm_reduce_mulsc_shrsc_sp33 & multm_reduce_mulsc_shrsc_cp33;
  assign multm_reduce_mulsc_shrsc_cq34 = multm_reduce_mulsc_shrsc_sp34 & multm_reduce_mulsc_shrsc_cp34;
  assign multm_reduce_mulsc_shrsc_cq35 = multm_reduce_mulsc_shrsc_sp35 & multm_reduce_mulsc_shrsc_cp35;
  assign multm_reduce_mulsc_shrsc_cq36 = multm_reduce_mulsc_shrsc_sp36 & multm_reduce_mulsc_shrsc_cp36;
  assign multm_reduce_mulsc_shrsc_cq37 = multm_reduce_mulsc_shrsc_sp37 & multm_reduce_mulsc_shrsc_cp37;
  assign multm_reduce_mulsc_shrsc_cq38 = multm_reduce_mulsc_shrsc_sp38 & multm_reduce_mulsc_shrsc_cp38;
  assign multm_reduce_mulsc_shrsc_cq39 = multm_reduce_mulsc_shrsc_sp39 & multm_reduce_mulsc_shrsc_cp39;
  assign multm_reduce_mulsc_shrsc_cq40 = multm_reduce_mulsc_shrsc_sp40 & multm_reduce_mulsc_shrsc_cp40;
  assign multm_reduce_mulsc_shrsc_cq41 = multm_reduce_mulsc_shrsc_sp41 & multm_reduce_mulsc_shrsc_cp41;
  assign multm_reduce_mulsc_shrsc_cq42 = multm_reduce_mulsc_shrsc_sp42 & multm_reduce_mulsc_shrsc_cp42;
  assign multm_reduce_mulsc_shrsc_cq43 = multm_reduce_mulsc_shrsc_sp43 & multm_reduce_mulsc_shrsc_cp43;
  assign multm_reduce_mulsc_shrsc_cq44 = multm_reduce_mulsc_shrsc_sp44 & multm_reduce_mulsc_shrsc_cp44;
  assign multm_reduce_mulsc_shrsc_cq45 = multm_reduce_mulsc_shrsc_sp45 & multm_reduce_mulsc_shrsc_cp45;
  assign multm_reduce_mulsc_shrsc_cq46 = multm_reduce_mulsc_shrsc_sp46 & multm_reduce_mulsc_shrsc_cp46;
  assign multm_reduce_mulsc_shrsc_cq47 = multm_reduce_mulsc_shrsc_sp47 & multm_reduce_mulsc_shrsc_cp47;
  assign multm_reduce_mulsc_shrsc_cq48 = multm_reduce_mulsc_shrsc_sp48 & multm_reduce_mulsc_shrsc_cp48;
  assign multm_reduce_mulsc_shrsc_cq49 = multm_reduce_mulsc_shrsc_sp49 & multm_reduce_mulsc_shrsc_cp49;
  assign multm_reduce_mulsc_shrsc_cq50 = multm_reduce_mulsc_shrsc_sp50 & multm_reduce_mulsc_shrsc_cp50;
  assign multm_reduce_mulsc_shrsc_cq51 = multm_reduce_mulsc_shrsc_sp51 & multm_reduce_mulsc_shrsc_cp51;
  assign multm_reduce_mulsc_shrsc_cq52 = multm_reduce_mulsc_shrsc_sp52 & multm_reduce_mulsc_shrsc_cp52;
  assign multm_reduce_mulsc_shrsc_cq53 = multm_reduce_mulsc_shrsc_sp53 & multm_reduce_mulsc_shrsc_cp53;
  assign multm_reduce_mulsc_shrsc_cq54 = multm_reduce_mulsc_shrsc_sp54 & multm_reduce_mulsc_shrsc_cp54;
  assign multm_reduce_mulsc_shrsc_cq55 = multm_reduce_mulsc_shrsc_sp55 & multm_reduce_mulsc_shrsc_cp55;
  assign multm_reduce_mulsc_shrsc_cq56 = multm_reduce_mulsc_shrsc_sp56 & multm_reduce_mulsc_shrsc_cp56;
  assign multm_reduce_mulsc_shrsc_cq57 = multm_reduce_mulsc_shrsc_sp57 & multm_reduce_mulsc_shrsc_cp57;
  assign multm_reduce_mulsc_shrsc_cq58 = multm_reduce_mulsc_shrsc_sp58 & multm_reduce_mulsc_shrsc_cp58;
  assign multm_reduce_mulsc_shrsc_cq59 = multm_reduce_mulsc_shrsc_sp59 & multm_reduce_mulsc_shrsc_cp59;
  assign multm_reduce_mulsc_shrsc_cq60 = multm_reduce_mulsc_shrsc_sp60 & multm_reduce_mulsc_shrsc_cp60;
  assign multm_reduce_mulsc_shrsc_cq61 = multm_reduce_mulsc_shrsc_sp61 & multm_reduce_mulsc_shrsc_cp61;
  assign multm_reduce_mulsc_shrsc_cq62 = multm_reduce_mulsc_shrsc_sp62 & multm_reduce_mulsc_shrsc_cp62;
  assign multm_reduce_mulsc_shrsc_cq63 = multm_reduce_mulsc_shrsc_sp63 & multm_reduce_mulsc_shrsc_cp63;
  assign multm_reduce_mulsc_shrsc_cq64 = multm_reduce_mulsc_shrsc_sp64 & multm_reduce_mulsc_shrsc_cp64;
  assign multm_reduce_mulsc_shrsc_cq65 = multm_reduce_mulsc_shrsc_sp65 & multm_reduce_mulsc_shrsc_cp65;
  assign multm_reduce_mulsc_shrsc_cq66 = multm_reduce_mulsc_shrsc_sp66 & multm_reduce_mulsc_shrsc_cp66;
  assign multm_reduce_mulsc_shrsc_cq67 = multm_reduce_mulsc_shrsc_sp67 & multm_reduce_mulsc_shrsc_cp67;
  assign multm_reduce_mulsc_shrsc_cq68 = multm_reduce_mulsc_shrsc_sp68 & multm_reduce_mulsc_shrsc_cp68;
  assign multm_reduce_mulsc_shrsc_cq69 = multm_reduce_mulsc_shrsc_sp69 & multm_reduce_mulsc_shrsc_cp69;
  assign multm_reduce_mulsc_shrsc_cq70 = multm_reduce_mulsc_shrsc_sp70 & multm_reduce_mulsc_shrsc_cp70;
  assign multm_reduce_mulsc_shrsc_cq71 = multm_reduce_mulsc_shrsc_sp71 & multm_reduce_mulsc_shrsc_cp71;
  assign multm_reduce_mulsc_shrsc_cq72 = multm_reduce_mulsc_shrsc_sp72 & multm_reduce_mulsc_shrsc_cp72;
  assign multm_reduce_mulsc_shrsc_cq73 = multm_reduce_mulsc_shrsc_sp73 & multm_reduce_mulsc_shrsc_cp73;
  assign multm_reduce_mulsc_shrsc_cq74 = multm_reduce_mulsc_shrsc_sp74 & multm_reduce_mulsc_shrsc_cp74;
  assign multm_reduce_mulsc_shrsc_cq75 = multm_reduce_mulsc_shrsc_sp75 & multm_reduce_mulsc_shrsc_cp75;
  assign multm_reduce_mulsc_shrsc_cq76 = multm_reduce_mulsc_shrsc_sp76 & multm_reduce_mulsc_shrsc_cp76;
  assign multm_reduce_mulsc_shrsc_cq77 = multm_reduce_mulsc_shrsc_sp77 & multm_reduce_mulsc_shrsc_cp77;
  assign multm_reduce_mulsc_shrsc_cq78 = multm_reduce_mulsc_shrsc_sp78 & multm_reduce_mulsc_shrsc_cp78;
  assign multm_reduce_mulsc_shrsc_cq79 = multm_reduce_mulsc_shrsc_sp79 & multm_reduce_mulsc_shrsc_cp79;
  assign multm_reduce_mulsc_shrsc_cq80 = multm_reduce_mulsc_shrsc_sp80 & multm_reduce_mulsc_shrsc_cp80;
  assign multm_reduce_mulsc_shrsc_cq81 = multm_reduce_mulsc_shrsc_sp81 & multm_reduce_mulsc_shrsc_cp81;
  assign multm_reduce_mulsc_shrsc_cq82 = multm_reduce_mulsc_shrsc_sp82 & multm_reduce_mulsc_shrsc_cp82;
  assign multm_reduce_mulsc_shrsc_cq83 = multm_reduce_mulsc_shrsc_sp83 & multm_reduce_mulsc_shrsc_cp83;
  assign multm_reduce_mulsc_shrsc_cq84 = multm_reduce_mulsc_shrsc_sp84 & multm_reduce_mulsc_shrsc_cp84;
  assign multm_reduce_mulsc_shrsc_cq85 = multm_reduce_mulsc_shrsc_sp85 & multm_reduce_mulsc_shrsc_cp85;
  assign multm_reduce_mulsc_shrsc_cq86 = multm_reduce_mulsc_shrsc_sp86 & multm_reduce_mulsc_shrsc_cp86;
  assign multm_reduce_mulsc_shrsc_cq87 = multm_reduce_mulsc_shrsc_sp87 & multm_reduce_mulsc_shrsc_cp87;
  assign multm_reduce_mulsc_shrsc_cq88 = multm_reduce_mulsc_shrsc_sp88 & multm_reduce_mulsc_shrsc_cp88;
  assign multm_reduce_mulsc_shrsc_cq89 = multm_reduce_mulsc_shrsc_sp89 & multm_reduce_mulsc_shrsc_cp89;
  assign multm_reduce_mulsc_shrsc_cq90 = multm_reduce_mulsc_shrsc_sp90 & multm_reduce_mulsc_shrsc_cp90;
  assign multm_reduce_mulsc_shrsc_cq91 = multm_reduce_mulsc_shrsc_sp91 & multm_reduce_mulsc_shrsc_cp91;
  assign multm_reduce_mulsc_shrsc_cq92 = multm_reduce_mulsc_shrsc_sp92 & multm_reduce_mulsc_shrsc_cp92;
  assign multm_reduce_mulsc_shrsc_cq93 = multm_reduce_mulsc_shrsc_sp93 & multm_reduce_mulsc_shrsc_cp93;
  assign multm_reduce_mulsc_shrsc_cq94 = multm_reduce_mulsc_shrsc_sp94 & multm_reduce_mulsc_shrsc_cp94;
  assign multm_reduce_mulsc_shrsc_cq95 = multm_reduce_mulsc_shrsc_sp95 & multm_reduce_mulsc_shrsc_cp95;
  assign multm_reduce_mulsc_shrsc_cq96 = multm_reduce_mulsc_shrsc_sp96 & multm_reduce_mulsc_shrsc_cp96;
  assign multm_reduce_mulsc_shrsc_cq97 = multm_reduce_mulsc_shrsc_sp97 & multm_reduce_mulsc_shrsc_cp97;
  assign multm_reduce_mulsc_shrsc_cq98 = multm_reduce_mulsc_shrsc_sp98 & multm_reduce_mulsc_shrsc_cp98;
  assign multm_reduce_mulsc_shrsc_cq99 = multm_reduce_mulsc_shrsc_sp99 & multm_reduce_mulsc_shrsc_cp99;
  assign multm_reduce_mulsc_shrsc_cq100 = multm_reduce_mulsc_shrsc_sp100 & multm_reduce_mulsc_shrsc_cp100;
  assign multm_reduce_mulsc_shrsc_cq101 = multm_reduce_mulsc_shrsc_sp101 & multm_reduce_mulsc_shrsc_cp101;
  assign multm_reduce_mulsc_shrsc_cq102 = multm_reduce_mulsc_shrsc_sp102 & multm_reduce_mulsc_shrsc_cp102;
  assign multm_reduce_mulsc_shrsc_cq103 = multm_reduce_mulsc_shrsc_sp103 & multm_reduce_mulsc_shrsc_cp103;
  assign multm_reduce_mulsc_shrsc_cq104 = multm_reduce_mulsc_shrsc_sp104 & multm_reduce_mulsc_shrsc_cp104;
  assign multm_reduce_mulsc_shrsc_cq105 = multm_reduce_mulsc_shrsc_sp105 & multm_reduce_mulsc_shrsc_cp105;
  assign multm_reduce_mulsc_shrsc_cq106 = multm_reduce_mulsc_shrsc_sp106 & multm_reduce_mulsc_shrsc_cp106;
  assign multm_reduce_mulsc_shrsc_cq107 = multm_reduce_mulsc_shrsc_sp107 & multm_reduce_mulsc_shrsc_cp107;
  assign multm_reduce_mulsc_shrsc_cq108 = multm_reduce_mulsc_shrsc_sp108 & multm_reduce_mulsc_shrsc_cp108;
  assign multm_reduce_mulsc_shrsc_cq109 = multm_reduce_mulsc_shrsc_sp109 & multm_reduce_mulsc_shrsc_cp109;
  assign multm_reduce_mulsc_shrsc_cq110 = multm_reduce_mulsc_shrsc_sp110 & multm_reduce_mulsc_shrsc_cp110;
  assign multm_reduce_mulsc_shrsc_cq111 = multm_reduce_mulsc_shrsc_sp111 & multm_reduce_mulsc_shrsc_cp111;
  assign multm_reduce_mulsc_shrsc_cq112 = multm_reduce_mulsc_shrsc_sp112 & multm_reduce_mulsc_shrsc_cp112;
  assign multm_reduce_mulsc_shrsc_cq113 = multm_reduce_mulsc_shrsc_sp113 & multm_reduce_mulsc_shrsc_cp113;
  assign multm_reduce_mulsc_shrsc_cq114 = multm_reduce_mulsc_shrsc_sp114 & multm_reduce_mulsc_shrsc_cp114;
  assign multm_reduce_mulsc_shrsc_cq115 = multm_reduce_mulsc_shrsc_sp115 & multm_reduce_mulsc_shrsc_cp115;
  assign multm_reduce_mulsc_shrsc_cq116 = multm_reduce_mulsc_shrsc_sp116 & multm_reduce_mulsc_shrsc_cp116;
  assign multm_reduce_mulsc_shrsc_cq117 = multm_reduce_mulsc_shrsc_sp117 & multm_reduce_mulsc_shrsc_cp117;
  assign multm_reduce_mulsc_shrsc_cq118 = multm_reduce_mulsc_shrsc_sp118 & multm_reduce_mulsc_shrsc_cp118;
  assign multm_reduce_mulsc_shrsc_cq119 = multm_reduce_mulsc_shrsc_sp119 & multm_reduce_mulsc_shrsc_cp119;
  assign multm_reduce_mulsc_shrsc_cq120 = multm_reduce_mulsc_shrsc_sp120 & multm_reduce_mulsc_shrsc_cp120;
  assign multm_reduce_mulsc_shrsc_cq121 = multm_reduce_mulsc_shrsc_sp121 & multm_reduce_mulsc_shrsc_cp121;
  assign multm_reduce_mulsc_shrsc_cq122 = multm_reduce_mulsc_shrsc_sp122 & multm_reduce_mulsc_shrsc_cp122;
  assign multm_reduce_mulsc_shrsc_cq123 = multm_reduce_mulsc_shrsc_sp123 & multm_reduce_mulsc_shrsc_cp123;
  assign multm_reduce_mulsc_shrsc_cq124 = multm_reduce_mulsc_shrsc_sp124 & multm_reduce_mulsc_shrsc_cp124;
  assign multm_reduce_mulsc_shrsc_cq125 = multm_reduce_mulsc_shrsc_sp125 & multm_reduce_mulsc_shrsc_cp125;
  assign multm_reduce_mulsc_shrsc_cq126 = multm_reduce_mulsc_shrsc_sp126 & multm_reduce_mulsc_shrsc_cp126;
  assign multm_reduce_mulsc_shrsc_cq127 = multm_reduce_mulsc_shrsc_sp127 & multm_reduce_mulsc_shrsc_cp127;
  assign multm_reduce_mulsc_shrsc_cq128 = multm_reduce_mulsc_shrsc_sp128 & multm_reduce_mulsc_shrsc_cp128;
  assign multm_reduce_mulsc_shrsc_cq129 = multm_reduce_mulsc_shrsc_sp129 & multm_reduce_mulsc_shrsc_cp129;
  assign multm_reduce_mulsc_shrsc_cq130 = multm_reduce_mulsc_shrsc_sp130 & multm_reduce_mulsc_shrsc_cp130;
  assign multm_reduce_mulsc_shrsc_cq131 = multm_reduce_mulsc_shrsc_sp131 & multm_reduce_mulsc_shrsc_cp131;
  assign multm_reduce_mulsc_shrsc_cq132 = multm_reduce_mulsc_shrsc_sp132 & multm_reduce_mulsc_shrsc_cp132;
  assign multm_reduce_mulsc_shrsc_cq133 = multm_reduce_mulsc_shrsc_sp133 & multm_reduce_mulsc_shrsc_cp133;
  assign multm_reduce_mulsc_shrsc_cq134 = multm_reduce_mulsc_shrsc_sp134 & multm_reduce_mulsc_shrsc_cp134;
  assign multm_reduce_mulsc_shrsc_cq135 = multm_reduce_mulsc_shrsc_sp135 & multm_reduce_mulsc_shrsc_cp135;
  assign multm_reduce_mulsc_shrsc_cq136 = multm_reduce_mulsc_shrsc_sp136 & multm_reduce_mulsc_shrsc_cp136;
  assign multm_reduce_mulsc_shrsc_cq137 = multm_reduce_mulsc_shrsc_sp137 & multm_reduce_mulsc_shrsc_cp137;
  assign multm_reduce_mulsc_shrsc_cq138 = multm_reduce_mulsc_shrsc_sp138 & multm_reduce_mulsc_shrsc_cp138;
  assign multm_reduce_mulsc_shrsc_cq139 = multm_reduce_mulsc_shrsc_sp139 & multm_reduce_mulsc_shrsc_cp139;
  assign multm_reduce_mulsc_shrsc_cq140 = multm_reduce_mulsc_shrsc_sp140 & multm_reduce_mulsc_shrsc_cp140;
  assign multm_reduce_mulsc_shrsc_cq141 = multm_reduce_mulsc_shrsc_sp141 & multm_reduce_mulsc_shrsc_cp141;
  assign multm_reduce_mulsc_shrsc_cq142 = multm_reduce_mulsc_shrsc_sp142 & multm_reduce_mulsc_shrsc_cp142;
  assign multm_reduce_mulsc_shrsc_cq143 = multm_reduce_mulsc_shrsc_sp143 & multm_reduce_mulsc_shrsc_cp143;
  assign multm_reduce_mulsc_shrsc_cq144 = multm_reduce_mulsc_shrsc_sp144 & multm_reduce_mulsc_shrsc_cp144;
  assign multm_reduce_mulsc_shrsc_cq145 = multm_reduce_mulsc_shrsc_sp145 & multm_reduce_mulsc_shrsc_cp145;
  assign multm_reduce_mulsc_shrsc_cq146 = multm_reduce_mulsc_shrsc_sp146 & multm_reduce_mulsc_shrsc_cp146;
  assign multm_reduce_mulsc_shrsc_cq147 = multm_reduce_mulsc_shrsc_sp147 & multm_reduce_mulsc_shrsc_cp147;
  assign multm_reduce_mulsc_shrsc_cq148 = multm_reduce_mulsc_shrsc_sp148 & multm_reduce_mulsc_shrsc_cp148;
  assign multm_reduce_mulsc_shrsc_cq149 = multm_reduce_mulsc_shrsc_sp149 & multm_reduce_mulsc_shrsc_cp149;
  assign multm_reduce_mulsc_shrsc_cq150 = multm_reduce_mulsc_shrsc_sp150 & multm_reduce_mulsc_shrsc_cp150;
  assign multm_reduce_mulsc_shrsc_cq151 = multm_reduce_mulsc_shrsc_sp151 & multm_reduce_mulsc_shrsc_cp151;
  assign multm_reduce_mulsc_shrsc_cq152 = multm_reduce_mulsc_shrsc_sp152 & multm_reduce_mulsc_shrsc_cp152;
  assign multm_reduce_mulsc_shrsc_cq153 = multm_reduce_mulsc_shrsc_sp153 & multm_reduce_mulsc_shrsc_cp153;
  assign multm_reduce_mulsc_shrsc_cq154 = multm_reduce_mulsc_shrsc_sp154 & multm_reduce_mulsc_shrsc_cp154;
  assign multm_reduce_mulsc_shrsc_cq155 = multm_reduce_mulsc_shrsc_sp155 & multm_reduce_mulsc_shrsc_cp155;
  assign multm_reduce_mulsc_shrsc_cq156 = multm_reduce_mulsc_shrsc_sp156 & multm_reduce_mulsc_shrsc_cp156;
  assign multm_reduce_mulsc_shrsc_cq157 = multm_reduce_mulsc_shrsc_sp157 & multm_reduce_mulsc_shrsc_cp157;
  assign multm_reduce_mulsc_shrsc_cq158 = multm_reduce_mulsc_shrsc_sp158 & multm_reduce_mulsc_shrsc_cp158;
  assign multm_reduce_mulsc_shrsc_cq159 = multm_reduce_mulsc_shrsc_sp159 & multm_reduce_mulsc_shrsc_cp159;
  assign multm_reduce_mulsc_shrsc_cq160 = multm_reduce_mulsc_shrsc_sp160 & multm_reduce_mulsc_shrsc_cp160;
  assign multm_reduce_mulsc_shrsc_cq161 = multm_reduce_mulsc_shrsc_sp161 & multm_reduce_mulsc_shrsc_cp161;
  assign multm_reduce_mulsc_shrsc_cq162 = multm_reduce_mulsc_shrsc_sp162 & multm_reduce_mulsc_shrsc_cp162;
  assign multm_reduce_mulsc_shrsc_cq163 = multm_reduce_mulsc_shrsc_sp163 & multm_reduce_mulsc_shrsc_cp163;
  assign multm_reduce_mulsc_shrsc_cq164 = multm_reduce_mulsc_shrsc_sp164 & multm_reduce_mulsc_shrsc_cp164;
  assign multm_reduce_mulsc_shrsc_cq165 = multm_reduce_mulsc_shrsc_sp165 & multm_reduce_mulsc_shrsc_cp165;
  assign multm_reduce_mulsc_shrsc_cq166 = multm_reduce_mulsc_shrsc_sp166 & multm_reduce_mulsc_shrsc_cp166;
  assign multm_reduce_mulsc_shrsc_cq167 = multm_reduce_mulsc_shrsc_sp167 & multm_reduce_mulsc_shrsc_cp167;
  assign multm_reduce_mulsc_shrsc_cq168 = multm_reduce_mulsc_shrsc_sp168 & multm_reduce_mulsc_shrsc_cp168;
  assign multm_reduce_mulsc_shrsc_cq169 = multm_reduce_mulsc_shrsc_sp169 & multm_reduce_mulsc_shrsc_cp169;
  assign multm_reduce_mulsc_shrsc_cq170 = multm_reduce_mulsc_shrsc_sp170 & multm_reduce_mulsc_shrsc_cp170;
  assign multm_reduce_mulsc_shrsc_cq171 = multm_reduce_mulsc_shrsc_sp171 & multm_reduce_mulsc_shrsc_cp171;
  assign multm_reduce_mulsc_shrsc_cq172 = multm_reduce_mulsc_shrsc_sp172 & multm_reduce_mulsc_shrsc_cp172;
  assign multm_reduce_mulsc_shrsc_cq173 = multm_reduce_mulsc_shrsc_sp173 & multm_reduce_mulsc_shrsc_cp173;
  assign multm_reduce_mulsc_shrsc_cq174 = multm_reduce_mulsc_shrsc_sp174 & multm_reduce_mulsc_shrsc_cp174;
  assign multm_reduce_mulsc_shrsc_cq175 = multm_reduce_mulsc_shrsc_sp175 & multm_reduce_mulsc_shrsc_cp175;
  assign multm_reduce_mulsc_shrsc_cq176 = multm_reduce_mulsc_shrsc_sp176 & multm_reduce_mulsc_shrsc_cp176;
  assign multm_reduce_mulsc_shrsc_cq177 = multm_reduce_mulsc_shrsc_sp177 & multm_reduce_mulsc_shrsc_cp177;
  assign multm_reduce_mulsc_shrsc_cq178 = multm_reduce_mulsc_shrsc_sp178 & multm_reduce_mulsc_shrsc_cp178;
  assign multm_reduce_mulsc_shrsc_cq179 = multm_reduce_mulsc_shrsc_sp179 & multm_reduce_mulsc_shrsc_cp179;
  assign multm_reduce_mulsc_shrsc_cq180 = multm_reduce_mulsc_shrsc_sp180 & multm_reduce_mulsc_shrsc_cp180;
  assign multm_reduce_mulsc_shrsc_cq181 = multm_reduce_mulsc_shrsc_sp181 & multm_reduce_mulsc_shrsc_cp181;
  assign multm_reduce_mulsc_shrsc_cq182 = multm_reduce_mulsc_shrsc_sp182 & multm_reduce_mulsc_shrsc_cp182;
  assign multm_reduce_mulsc_shrsc_cr0 = sadd ? yc0_o : multm_reduce_mulsc_shrsc_cq0;
  assign multm_reduce_mulsc_shrsc_cr1 = sadd ? yc1_o : multm_reduce_mulsc_shrsc_cq1;
  assign multm_reduce_mulsc_shrsc_cr2 = sadd ? yc2_o : multm_reduce_mulsc_shrsc_cq2;
  assign multm_reduce_mulsc_shrsc_cr3 = sadd ? yc3_o : multm_reduce_mulsc_shrsc_cq3;
  assign multm_reduce_mulsc_shrsc_cr4 = sadd ? yc4_o : multm_reduce_mulsc_shrsc_cq4;
  assign multm_reduce_mulsc_shrsc_cr5 = sadd ? yc5_o : multm_reduce_mulsc_shrsc_cq5;
  assign multm_reduce_mulsc_shrsc_cr6 = sadd ? yc6_o : multm_reduce_mulsc_shrsc_cq6;
  assign multm_reduce_mulsc_shrsc_cr7 = sadd ? yc7_o : multm_reduce_mulsc_shrsc_cq7;
  assign multm_reduce_mulsc_shrsc_cr8 = sadd ? yc8_o : multm_reduce_mulsc_shrsc_cq8;
  assign multm_reduce_mulsc_shrsc_cr9 = sadd ? yc9_o : multm_reduce_mulsc_shrsc_cq9;
  assign multm_reduce_mulsc_shrsc_cr10 = sadd ? yc10_o : multm_reduce_mulsc_shrsc_cq10;
  assign multm_reduce_mulsc_shrsc_cr11 = sadd ? yc11_o : multm_reduce_mulsc_shrsc_cq11;
  assign multm_reduce_mulsc_shrsc_cr12 = sadd ? yc12_o : multm_reduce_mulsc_shrsc_cq12;
  assign multm_reduce_mulsc_shrsc_cr13 = sadd ? yc13_o : multm_reduce_mulsc_shrsc_cq13;
  assign multm_reduce_mulsc_shrsc_cr14 = sadd ? yc14_o : multm_reduce_mulsc_shrsc_cq14;
  assign multm_reduce_mulsc_shrsc_cr15 = sadd ? yc15_o : multm_reduce_mulsc_shrsc_cq15;
  assign multm_reduce_mulsc_shrsc_cr16 = sadd ? yc16_o : multm_reduce_mulsc_shrsc_cq16;
  assign multm_reduce_mulsc_shrsc_cr17 = sadd ? yc17_o : multm_reduce_mulsc_shrsc_cq17;
  assign multm_reduce_mulsc_shrsc_cr18 = sadd ? yc18_o : multm_reduce_mulsc_shrsc_cq18;
  assign multm_reduce_mulsc_shrsc_cr19 = sadd ? yc19_o : multm_reduce_mulsc_shrsc_cq19;
  assign multm_reduce_mulsc_shrsc_cr20 = sadd ? yc20_o : multm_reduce_mulsc_shrsc_cq20;
  assign multm_reduce_mulsc_shrsc_cr21 = sadd ? yc21_o : multm_reduce_mulsc_shrsc_cq21;
  assign multm_reduce_mulsc_shrsc_cr22 = sadd ? yc22_o : multm_reduce_mulsc_shrsc_cq22;
  assign multm_reduce_mulsc_shrsc_cr23 = sadd ? yc23_o : multm_reduce_mulsc_shrsc_cq23;
  assign multm_reduce_mulsc_shrsc_cr24 = sadd ? yc24_o : multm_reduce_mulsc_shrsc_cq24;
  assign multm_reduce_mulsc_shrsc_cr25 = sadd ? yc25_o : multm_reduce_mulsc_shrsc_cq25;
  assign multm_reduce_mulsc_shrsc_cr26 = sadd ? yc26_o : multm_reduce_mulsc_shrsc_cq26;
  assign multm_reduce_mulsc_shrsc_cr27 = sadd ? yc27_o : multm_reduce_mulsc_shrsc_cq27;
  assign multm_reduce_mulsc_shrsc_cr28 = sadd ? yc28_o : multm_reduce_mulsc_shrsc_cq28;
  assign multm_reduce_mulsc_shrsc_cr29 = sadd ? yc29_o : multm_reduce_mulsc_shrsc_cq29;
  assign multm_reduce_mulsc_shrsc_cr30 = sadd ? yc30_o : multm_reduce_mulsc_shrsc_cq30;
  assign multm_reduce_mulsc_shrsc_cr31 = sadd ? yc31_o : multm_reduce_mulsc_shrsc_cq31;
  assign multm_reduce_mulsc_shrsc_cr32 = sadd ? yc32_o : multm_reduce_mulsc_shrsc_cq32;
  assign multm_reduce_mulsc_shrsc_cr33 = sadd ? yc33_o : multm_reduce_mulsc_shrsc_cq33;
  assign multm_reduce_mulsc_shrsc_cr34 = sadd ? yc34_o : multm_reduce_mulsc_shrsc_cq34;
  assign multm_reduce_mulsc_shrsc_cr35 = sadd ? yc35_o : multm_reduce_mulsc_shrsc_cq35;
  assign multm_reduce_mulsc_shrsc_cr36 = sadd ? yc36_o : multm_reduce_mulsc_shrsc_cq36;
  assign multm_reduce_mulsc_shrsc_cr37 = sadd ? yc37_o : multm_reduce_mulsc_shrsc_cq37;
  assign multm_reduce_mulsc_shrsc_cr38 = sadd ? yc38_o : multm_reduce_mulsc_shrsc_cq38;
  assign multm_reduce_mulsc_shrsc_cr39 = sadd ? yc39_o : multm_reduce_mulsc_shrsc_cq39;
  assign multm_reduce_mulsc_shrsc_cr40 = sadd ? yc40_o : multm_reduce_mulsc_shrsc_cq40;
  assign multm_reduce_mulsc_shrsc_cr41 = sadd ? yc41_o : multm_reduce_mulsc_shrsc_cq41;
  assign multm_reduce_mulsc_shrsc_cr42 = sadd ? yc42_o : multm_reduce_mulsc_shrsc_cq42;
  assign multm_reduce_mulsc_shrsc_cr43 = sadd ? yc43_o : multm_reduce_mulsc_shrsc_cq43;
  assign multm_reduce_mulsc_shrsc_cr44 = sadd ? yc44_o : multm_reduce_mulsc_shrsc_cq44;
  assign multm_reduce_mulsc_shrsc_cr45 = sadd ? yc45_o : multm_reduce_mulsc_shrsc_cq45;
  assign multm_reduce_mulsc_shrsc_cr46 = sadd ? yc46_o : multm_reduce_mulsc_shrsc_cq46;
  assign multm_reduce_mulsc_shrsc_cr47 = sadd ? yc47_o : multm_reduce_mulsc_shrsc_cq47;
  assign multm_reduce_mulsc_shrsc_cr48 = sadd ? yc48_o : multm_reduce_mulsc_shrsc_cq48;
  assign multm_reduce_mulsc_shrsc_cr49 = sadd ? yc49_o : multm_reduce_mulsc_shrsc_cq49;
  assign multm_reduce_mulsc_shrsc_cr50 = sadd ? yc50_o : multm_reduce_mulsc_shrsc_cq50;
  assign multm_reduce_mulsc_shrsc_cr51 = sadd ? yc51_o : multm_reduce_mulsc_shrsc_cq51;
  assign multm_reduce_mulsc_shrsc_cr52 = sadd ? yc52_o : multm_reduce_mulsc_shrsc_cq52;
  assign multm_reduce_mulsc_shrsc_cr53 = sadd ? yc53_o : multm_reduce_mulsc_shrsc_cq53;
  assign multm_reduce_mulsc_shrsc_cr54 = sadd ? yc54_o : multm_reduce_mulsc_shrsc_cq54;
  assign multm_reduce_mulsc_shrsc_cr55 = sadd ? yc55_o : multm_reduce_mulsc_shrsc_cq55;
  assign multm_reduce_mulsc_shrsc_cr56 = sadd ? yc56_o : multm_reduce_mulsc_shrsc_cq56;
  assign multm_reduce_mulsc_shrsc_cr57 = sadd ? yc57_o : multm_reduce_mulsc_shrsc_cq57;
  assign multm_reduce_mulsc_shrsc_cr58 = sadd ? yc58_o : multm_reduce_mulsc_shrsc_cq58;
  assign multm_reduce_mulsc_shrsc_cr59 = sadd ? yc59_o : multm_reduce_mulsc_shrsc_cq59;
  assign multm_reduce_mulsc_shrsc_cr60 = sadd ? yc60_o : multm_reduce_mulsc_shrsc_cq60;
  assign multm_reduce_mulsc_shrsc_cr61 = sadd ? yc61_o : multm_reduce_mulsc_shrsc_cq61;
  assign multm_reduce_mulsc_shrsc_cr62 = sadd ? yc62_o : multm_reduce_mulsc_shrsc_cq62;
  assign multm_reduce_mulsc_shrsc_cr63 = sadd ? yc63_o : multm_reduce_mulsc_shrsc_cq63;
  assign multm_reduce_mulsc_shrsc_cr64 = sadd ? yc64_o : multm_reduce_mulsc_shrsc_cq64;
  assign multm_reduce_mulsc_shrsc_cr65 = sadd ? yc65_o : multm_reduce_mulsc_shrsc_cq65;
  assign multm_reduce_mulsc_shrsc_cr66 = sadd ? yc66_o : multm_reduce_mulsc_shrsc_cq66;
  assign multm_reduce_mulsc_shrsc_cr67 = sadd ? yc67_o : multm_reduce_mulsc_shrsc_cq67;
  assign multm_reduce_mulsc_shrsc_cr68 = sadd ? yc68_o : multm_reduce_mulsc_shrsc_cq68;
  assign multm_reduce_mulsc_shrsc_cr69 = sadd ? yc69_o : multm_reduce_mulsc_shrsc_cq69;
  assign multm_reduce_mulsc_shrsc_cr70 = sadd ? yc70_o : multm_reduce_mulsc_shrsc_cq70;
  assign multm_reduce_mulsc_shrsc_cr71 = sadd ? yc71_o : multm_reduce_mulsc_shrsc_cq71;
  assign multm_reduce_mulsc_shrsc_cr72 = sadd ? yc72_o : multm_reduce_mulsc_shrsc_cq72;
  assign multm_reduce_mulsc_shrsc_cr73 = sadd ? yc73_o : multm_reduce_mulsc_shrsc_cq73;
  assign multm_reduce_mulsc_shrsc_cr74 = sadd ? yc74_o : multm_reduce_mulsc_shrsc_cq74;
  assign multm_reduce_mulsc_shrsc_cr75 = sadd ? yc75_o : multm_reduce_mulsc_shrsc_cq75;
  assign multm_reduce_mulsc_shrsc_cr76 = sadd ? yc76_o : multm_reduce_mulsc_shrsc_cq76;
  assign multm_reduce_mulsc_shrsc_cr77 = sadd ? yc77_o : multm_reduce_mulsc_shrsc_cq77;
  assign multm_reduce_mulsc_shrsc_cr78 = sadd ? yc78_o : multm_reduce_mulsc_shrsc_cq78;
  assign multm_reduce_mulsc_shrsc_cr79 = sadd ? yc79_o : multm_reduce_mulsc_shrsc_cq79;
  assign multm_reduce_mulsc_shrsc_cr80 = sadd ? yc80_o : multm_reduce_mulsc_shrsc_cq80;
  assign multm_reduce_mulsc_shrsc_cr81 = sadd ? yc81_o : multm_reduce_mulsc_shrsc_cq81;
  assign multm_reduce_mulsc_shrsc_cr82 = sadd ? yc82_o : multm_reduce_mulsc_shrsc_cq82;
  assign multm_reduce_mulsc_shrsc_cr83 = sadd ? yc83_o : multm_reduce_mulsc_shrsc_cq83;
  assign multm_reduce_mulsc_shrsc_cr84 = sadd ? yc84_o : multm_reduce_mulsc_shrsc_cq84;
  assign multm_reduce_mulsc_shrsc_cr85 = sadd ? yc85_o : multm_reduce_mulsc_shrsc_cq85;
  assign multm_reduce_mulsc_shrsc_cr86 = sadd ? yc86_o : multm_reduce_mulsc_shrsc_cq86;
  assign multm_reduce_mulsc_shrsc_cr87 = sadd ? yc87_o : multm_reduce_mulsc_shrsc_cq87;
  assign multm_reduce_mulsc_shrsc_cr88 = sadd ? yc88_o : multm_reduce_mulsc_shrsc_cq88;
  assign multm_reduce_mulsc_shrsc_cr89 = sadd ? yc89_o : multm_reduce_mulsc_shrsc_cq89;
  assign multm_reduce_mulsc_shrsc_cr90 = sadd ? yc90_o : multm_reduce_mulsc_shrsc_cq90;
  assign multm_reduce_mulsc_shrsc_cr91 = sadd ? yc91_o : multm_reduce_mulsc_shrsc_cq91;
  assign multm_reduce_mulsc_shrsc_cr92 = sadd ? yc92_o : multm_reduce_mulsc_shrsc_cq92;
  assign multm_reduce_mulsc_shrsc_cr93 = sadd ? yc93_o : multm_reduce_mulsc_shrsc_cq93;
  assign multm_reduce_mulsc_shrsc_cr94 = sadd ? yc94_o : multm_reduce_mulsc_shrsc_cq94;
  assign multm_reduce_mulsc_shrsc_cr95 = sadd ? yc95_o : multm_reduce_mulsc_shrsc_cq95;
  assign multm_reduce_mulsc_shrsc_cr96 = sadd ? yc96_o : multm_reduce_mulsc_shrsc_cq96;
  assign multm_reduce_mulsc_shrsc_cr97 = sadd ? yc97_o : multm_reduce_mulsc_shrsc_cq97;
  assign multm_reduce_mulsc_shrsc_cr98 = sadd ? yc98_o : multm_reduce_mulsc_shrsc_cq98;
  assign multm_reduce_mulsc_shrsc_cr99 = sadd ? yc99_o : multm_reduce_mulsc_shrsc_cq99;
  assign multm_reduce_mulsc_shrsc_cr100 = sadd ? yc100_o : multm_reduce_mulsc_shrsc_cq100;
  assign multm_reduce_mulsc_shrsc_cr101 = sadd ? yc101_o : multm_reduce_mulsc_shrsc_cq101;
  assign multm_reduce_mulsc_shrsc_cr102 = sadd ? yc102_o : multm_reduce_mulsc_shrsc_cq102;
  assign multm_reduce_mulsc_shrsc_cr103 = sadd ? yc103_o : multm_reduce_mulsc_shrsc_cq103;
  assign multm_reduce_mulsc_shrsc_cr104 = sadd ? yc104_o : multm_reduce_mulsc_shrsc_cq104;
  assign multm_reduce_mulsc_shrsc_cr105 = sadd ? yc105_o : multm_reduce_mulsc_shrsc_cq105;
  assign multm_reduce_mulsc_shrsc_cr106 = sadd ? yc106_o : multm_reduce_mulsc_shrsc_cq106;
  assign multm_reduce_mulsc_shrsc_cr107 = sadd ? yc107_o : multm_reduce_mulsc_shrsc_cq107;
  assign multm_reduce_mulsc_shrsc_cr108 = sadd ? yc108_o : multm_reduce_mulsc_shrsc_cq108;
  assign multm_reduce_mulsc_shrsc_cr109 = sadd ? yc109_o : multm_reduce_mulsc_shrsc_cq109;
  assign multm_reduce_mulsc_shrsc_cr110 = sadd ? yc110_o : multm_reduce_mulsc_shrsc_cq110;
  assign multm_reduce_mulsc_shrsc_cr111 = sadd ? yc111_o : multm_reduce_mulsc_shrsc_cq111;
  assign multm_reduce_mulsc_shrsc_cr112 = sadd ? yc112_o : multm_reduce_mulsc_shrsc_cq112;
  assign multm_reduce_mulsc_shrsc_cr113 = sadd ? yc113_o : multm_reduce_mulsc_shrsc_cq113;
  assign multm_reduce_mulsc_shrsc_cr114 = sadd ? yc114_o : multm_reduce_mulsc_shrsc_cq114;
  assign multm_reduce_mulsc_shrsc_cr115 = sadd ? yc115_o : multm_reduce_mulsc_shrsc_cq115;
  assign multm_reduce_mulsc_shrsc_cr116 = sadd ? yc116_o : multm_reduce_mulsc_shrsc_cq116;
  assign multm_reduce_mulsc_shrsc_cr117 = sadd ? yc117_o : multm_reduce_mulsc_shrsc_cq117;
  assign multm_reduce_mulsc_shrsc_cr118 = sadd ? yc118_o : multm_reduce_mulsc_shrsc_cq118;
  assign multm_reduce_mulsc_shrsc_cr119 = sadd ? yc119_o : multm_reduce_mulsc_shrsc_cq119;
  assign multm_reduce_mulsc_shrsc_cr120 = sadd ? yc120_o : multm_reduce_mulsc_shrsc_cq120;
  assign multm_reduce_mulsc_shrsc_cr121 = sadd ? yc121_o : multm_reduce_mulsc_shrsc_cq121;
  assign multm_reduce_mulsc_shrsc_cr122 = sadd ? yc122_o : multm_reduce_mulsc_shrsc_cq122;
  assign multm_reduce_mulsc_shrsc_cr123 = sadd ? yc123_o : multm_reduce_mulsc_shrsc_cq123;
  assign multm_reduce_mulsc_shrsc_cr124 = sadd ? yc124_o : multm_reduce_mulsc_shrsc_cq124;
  assign multm_reduce_mulsc_shrsc_cr125 = sadd ? yc125_o : multm_reduce_mulsc_shrsc_cq125;
  assign multm_reduce_mulsc_shrsc_cr126 = sadd ? yc126_o : multm_reduce_mulsc_shrsc_cq126;
  assign multm_reduce_mulsc_shrsc_cr127 = sadd ? yc127_o : multm_reduce_mulsc_shrsc_cq127;
  assign multm_reduce_mulsc_shrsc_cr128 = sadd ? yc128_o : multm_reduce_mulsc_shrsc_cq128;
  assign multm_reduce_mulsc_shrsc_cr129 = sadd ? yc129_o : multm_reduce_mulsc_shrsc_cq129;
  assign multm_reduce_mulsc_shrsc_cr130 = sadd ? yc130_o : multm_reduce_mulsc_shrsc_cq130;
  assign multm_reduce_mulsc_shrsc_cr131 = sadd ? yc131_o : multm_reduce_mulsc_shrsc_cq131;
  assign multm_reduce_mulsc_shrsc_cr132 = sadd ? yc132_o : multm_reduce_mulsc_shrsc_cq132;
  assign multm_reduce_mulsc_shrsc_cr133 = sadd ? yc133_o : multm_reduce_mulsc_shrsc_cq133;
  assign multm_reduce_mulsc_shrsc_cr134 = sadd ? yc134_o : multm_reduce_mulsc_shrsc_cq134;
  assign multm_reduce_mulsc_shrsc_cr135 = sadd ? yc135_o : multm_reduce_mulsc_shrsc_cq135;
  assign multm_reduce_mulsc_shrsc_cr136 = sadd ? yc136_o : multm_reduce_mulsc_shrsc_cq136;
  assign multm_reduce_mulsc_shrsc_cr137 = sadd ? yc137_o : multm_reduce_mulsc_shrsc_cq137;
  assign multm_reduce_mulsc_shrsc_cr138 = sadd ? yc138_o : multm_reduce_mulsc_shrsc_cq138;
  assign multm_reduce_mulsc_shrsc_cr139 = sadd ? yc139_o : multm_reduce_mulsc_shrsc_cq139;
  assign multm_reduce_mulsc_shrsc_cr140 = sadd ? yc140_o : multm_reduce_mulsc_shrsc_cq140;
  assign multm_reduce_mulsc_shrsc_cr141 = sadd ? yc141_o : multm_reduce_mulsc_shrsc_cq141;
  assign multm_reduce_mulsc_shrsc_cr142 = sadd ? yc142_o : multm_reduce_mulsc_shrsc_cq142;
  assign multm_reduce_mulsc_shrsc_cr143 = sadd ? yc143_o : multm_reduce_mulsc_shrsc_cq143;
  assign multm_reduce_mulsc_shrsc_cr144 = sadd ? yc144_o : multm_reduce_mulsc_shrsc_cq144;
  assign multm_reduce_mulsc_shrsc_cr145 = sadd ? yc145_o : multm_reduce_mulsc_shrsc_cq145;
  assign multm_reduce_mulsc_shrsc_cr146 = sadd ? yc146_o : multm_reduce_mulsc_shrsc_cq146;
  assign multm_reduce_mulsc_shrsc_cr147 = sadd ? yc147_o : multm_reduce_mulsc_shrsc_cq147;
  assign multm_reduce_mulsc_shrsc_cr148 = sadd ? yc148_o : multm_reduce_mulsc_shrsc_cq148;
  assign multm_reduce_mulsc_shrsc_cr149 = sadd ? yc149_o : multm_reduce_mulsc_shrsc_cq149;
  assign multm_reduce_mulsc_shrsc_cr150 = sadd ? yc150_o : multm_reduce_mulsc_shrsc_cq150;
  assign multm_reduce_mulsc_shrsc_cr151 = sadd ? yc151_o : multm_reduce_mulsc_shrsc_cq151;
  assign multm_reduce_mulsc_shrsc_cr152 = sadd ? yc152_o : multm_reduce_mulsc_shrsc_cq152;
  assign multm_reduce_mulsc_shrsc_cr153 = sadd ? yc153_o : multm_reduce_mulsc_shrsc_cq153;
  assign multm_reduce_mulsc_shrsc_cr154 = sadd ? yc154_o : multm_reduce_mulsc_shrsc_cq154;
  assign multm_reduce_mulsc_shrsc_cr155 = sadd ? yc155_o : multm_reduce_mulsc_shrsc_cq155;
  assign multm_reduce_mulsc_shrsc_cr156 = sadd ? yc156_o : multm_reduce_mulsc_shrsc_cq156;
  assign multm_reduce_mulsc_shrsc_cr157 = sadd ? yc157_o : multm_reduce_mulsc_shrsc_cq157;
  assign multm_reduce_mulsc_shrsc_cr158 = sadd ? yc158_o : multm_reduce_mulsc_shrsc_cq158;
  assign multm_reduce_mulsc_shrsc_cr159 = sadd ? yc159_o : multm_reduce_mulsc_shrsc_cq159;
  assign multm_reduce_mulsc_shrsc_cr160 = sadd ? yc160_o : multm_reduce_mulsc_shrsc_cq160;
  assign multm_reduce_mulsc_shrsc_cr161 = sadd ? yc161_o : multm_reduce_mulsc_shrsc_cq161;
  assign multm_reduce_mulsc_shrsc_cr162 = sadd ? yc162_o : multm_reduce_mulsc_shrsc_cq162;
  assign multm_reduce_mulsc_shrsc_cr163 = sadd ? yc163_o : multm_reduce_mulsc_shrsc_cq163;
  assign multm_reduce_mulsc_shrsc_cr164 = sadd ? yc164_o : multm_reduce_mulsc_shrsc_cq164;
  assign multm_reduce_mulsc_shrsc_cr165 = sadd ? yc165_o : multm_reduce_mulsc_shrsc_cq165;
  assign multm_reduce_mulsc_shrsc_cr166 = sadd ? yc166_o : multm_reduce_mulsc_shrsc_cq166;
  assign multm_reduce_mulsc_shrsc_cr167 = sadd ? yc167_o : multm_reduce_mulsc_shrsc_cq167;
  assign multm_reduce_mulsc_shrsc_cr168 = sadd ? yc168_o : multm_reduce_mulsc_shrsc_cq168;
  assign multm_reduce_mulsc_shrsc_cr169 = sadd ? yc169_o : multm_reduce_mulsc_shrsc_cq169;
  assign multm_reduce_mulsc_shrsc_cr170 = sadd ? yc170_o : multm_reduce_mulsc_shrsc_cq170;
  assign multm_reduce_mulsc_shrsc_cr171 = sadd ? yc171_o : multm_reduce_mulsc_shrsc_cq171;
  assign multm_reduce_mulsc_shrsc_cr172 = sadd ? yc172_o : multm_reduce_mulsc_shrsc_cq172;
  assign multm_reduce_mulsc_shrsc_cr173 = sadd ? yc173_o : multm_reduce_mulsc_shrsc_cq173;
  assign multm_reduce_mulsc_shrsc_cr174 = sadd ? yc174_o : multm_reduce_mulsc_shrsc_cq174;
  assign multm_reduce_mulsc_shrsc_cr175 = sadd ? yc175_o : multm_reduce_mulsc_shrsc_cq175;
  assign multm_reduce_mulsc_shrsc_cr176 = sadd ? yc176_o : multm_reduce_mulsc_shrsc_cq176;
  assign multm_reduce_mulsc_shrsc_cr177 = sadd ? yc177_o : multm_reduce_mulsc_shrsc_cq177;
  assign multm_reduce_mulsc_shrsc_cr178 = sadd ? yc178_o : multm_reduce_mulsc_shrsc_cq178;
  assign multm_reduce_mulsc_shrsc_cr179 = sadd ? yc179_o : multm_reduce_mulsc_shrsc_cq179;
  assign multm_reduce_mulsc_shrsc_cr180 = sadd ? yc180_o : multm_reduce_mulsc_shrsc_cq180;
  assign multm_reduce_mulsc_shrsc_cr181 = sadd ? yc181_o : multm_reduce_mulsc_shrsc_cq181;
  assign multm_reduce_mulsc_shrsc_cr182 = sadd ? yc182_o : multm_reduce_mulsc_shrsc_cq182;
  assign multm_reduce_mulsc_shrsc_cr183 = sadd & yc183_o;
  assign multm_reduce_mulsc_shrsc_sq0 = multm_reduce_mulsc_shrsc_sp0 ^ multm_reduce_mulsc_shrsc_cp0;
  assign multm_reduce_mulsc_shrsc_sq1 = multm_reduce_mulsc_shrsc_sp1 ^ multm_reduce_mulsc_shrsc_cp1;
  assign multm_reduce_mulsc_shrsc_sq2 = multm_reduce_mulsc_shrsc_sp2 ^ multm_reduce_mulsc_shrsc_cp2;
  assign multm_reduce_mulsc_shrsc_sq3 = multm_reduce_mulsc_shrsc_sp3 ^ multm_reduce_mulsc_shrsc_cp3;
  assign multm_reduce_mulsc_shrsc_sq4 = multm_reduce_mulsc_shrsc_sp4 ^ multm_reduce_mulsc_shrsc_cp4;
  assign multm_reduce_mulsc_shrsc_sq5 = multm_reduce_mulsc_shrsc_sp5 ^ multm_reduce_mulsc_shrsc_cp5;
  assign multm_reduce_mulsc_shrsc_sq6 = multm_reduce_mulsc_shrsc_sp6 ^ multm_reduce_mulsc_shrsc_cp6;
  assign multm_reduce_mulsc_shrsc_sq7 = multm_reduce_mulsc_shrsc_sp7 ^ multm_reduce_mulsc_shrsc_cp7;
  assign multm_reduce_mulsc_shrsc_sq8 = multm_reduce_mulsc_shrsc_sp8 ^ multm_reduce_mulsc_shrsc_cp8;
  assign multm_reduce_mulsc_shrsc_sq9 = multm_reduce_mulsc_shrsc_sp9 ^ multm_reduce_mulsc_shrsc_cp9;
  assign multm_reduce_mulsc_shrsc_sq10 = multm_reduce_mulsc_shrsc_sp10 ^ multm_reduce_mulsc_shrsc_cp10;
  assign multm_reduce_mulsc_shrsc_sq11 = multm_reduce_mulsc_shrsc_sp11 ^ multm_reduce_mulsc_shrsc_cp11;
  assign multm_reduce_mulsc_shrsc_sq12 = multm_reduce_mulsc_shrsc_sp12 ^ multm_reduce_mulsc_shrsc_cp12;
  assign multm_reduce_mulsc_shrsc_sq13 = multm_reduce_mulsc_shrsc_sp13 ^ multm_reduce_mulsc_shrsc_cp13;
  assign multm_reduce_mulsc_shrsc_sq14 = multm_reduce_mulsc_shrsc_sp14 ^ multm_reduce_mulsc_shrsc_cp14;
  assign multm_reduce_mulsc_shrsc_sq15 = multm_reduce_mulsc_shrsc_sp15 ^ multm_reduce_mulsc_shrsc_cp15;
  assign multm_reduce_mulsc_shrsc_sq16 = multm_reduce_mulsc_shrsc_sp16 ^ multm_reduce_mulsc_shrsc_cp16;
  assign multm_reduce_mulsc_shrsc_sq17 = multm_reduce_mulsc_shrsc_sp17 ^ multm_reduce_mulsc_shrsc_cp17;
  assign multm_reduce_mulsc_shrsc_sq18 = multm_reduce_mulsc_shrsc_sp18 ^ multm_reduce_mulsc_shrsc_cp18;
  assign multm_reduce_mulsc_shrsc_sq19 = multm_reduce_mulsc_shrsc_sp19 ^ multm_reduce_mulsc_shrsc_cp19;
  assign multm_reduce_mulsc_shrsc_sq20 = multm_reduce_mulsc_shrsc_sp20 ^ multm_reduce_mulsc_shrsc_cp20;
  assign multm_reduce_mulsc_shrsc_sq21 = multm_reduce_mulsc_shrsc_sp21 ^ multm_reduce_mulsc_shrsc_cp21;
  assign multm_reduce_mulsc_shrsc_sq22 = multm_reduce_mulsc_shrsc_sp22 ^ multm_reduce_mulsc_shrsc_cp22;
  assign multm_reduce_mulsc_shrsc_sq23 = multm_reduce_mulsc_shrsc_sp23 ^ multm_reduce_mulsc_shrsc_cp23;
  assign multm_reduce_mulsc_shrsc_sq24 = multm_reduce_mulsc_shrsc_sp24 ^ multm_reduce_mulsc_shrsc_cp24;
  assign multm_reduce_mulsc_shrsc_sq25 = multm_reduce_mulsc_shrsc_sp25 ^ multm_reduce_mulsc_shrsc_cp25;
  assign multm_reduce_mulsc_shrsc_sq26 = multm_reduce_mulsc_shrsc_sp26 ^ multm_reduce_mulsc_shrsc_cp26;
  assign multm_reduce_mulsc_shrsc_sq27 = multm_reduce_mulsc_shrsc_sp27 ^ multm_reduce_mulsc_shrsc_cp27;
  assign multm_reduce_mulsc_shrsc_sq28 = multm_reduce_mulsc_shrsc_sp28 ^ multm_reduce_mulsc_shrsc_cp28;
  assign multm_reduce_mulsc_shrsc_sq29 = multm_reduce_mulsc_shrsc_sp29 ^ multm_reduce_mulsc_shrsc_cp29;
  assign multm_reduce_mulsc_shrsc_sq30 = multm_reduce_mulsc_shrsc_sp30 ^ multm_reduce_mulsc_shrsc_cp30;
  assign multm_reduce_mulsc_shrsc_sq31 = multm_reduce_mulsc_shrsc_sp31 ^ multm_reduce_mulsc_shrsc_cp31;
  assign multm_reduce_mulsc_shrsc_sq32 = multm_reduce_mulsc_shrsc_sp32 ^ multm_reduce_mulsc_shrsc_cp32;
  assign multm_reduce_mulsc_shrsc_sq33 = multm_reduce_mulsc_shrsc_sp33 ^ multm_reduce_mulsc_shrsc_cp33;
  assign multm_reduce_mulsc_shrsc_sq34 = multm_reduce_mulsc_shrsc_sp34 ^ multm_reduce_mulsc_shrsc_cp34;
  assign multm_reduce_mulsc_shrsc_sq35 = multm_reduce_mulsc_shrsc_sp35 ^ multm_reduce_mulsc_shrsc_cp35;
  assign multm_reduce_mulsc_shrsc_sq36 = multm_reduce_mulsc_shrsc_sp36 ^ multm_reduce_mulsc_shrsc_cp36;
  assign multm_reduce_mulsc_shrsc_sq37 = multm_reduce_mulsc_shrsc_sp37 ^ multm_reduce_mulsc_shrsc_cp37;
  assign multm_reduce_mulsc_shrsc_sq38 = multm_reduce_mulsc_shrsc_sp38 ^ multm_reduce_mulsc_shrsc_cp38;
  assign multm_reduce_mulsc_shrsc_sq39 = multm_reduce_mulsc_shrsc_sp39 ^ multm_reduce_mulsc_shrsc_cp39;
  assign multm_reduce_mulsc_shrsc_sq40 = multm_reduce_mulsc_shrsc_sp40 ^ multm_reduce_mulsc_shrsc_cp40;
  assign multm_reduce_mulsc_shrsc_sq41 = multm_reduce_mulsc_shrsc_sp41 ^ multm_reduce_mulsc_shrsc_cp41;
  assign multm_reduce_mulsc_shrsc_sq42 = multm_reduce_mulsc_shrsc_sp42 ^ multm_reduce_mulsc_shrsc_cp42;
  assign multm_reduce_mulsc_shrsc_sq43 = multm_reduce_mulsc_shrsc_sp43 ^ multm_reduce_mulsc_shrsc_cp43;
  assign multm_reduce_mulsc_shrsc_sq44 = multm_reduce_mulsc_shrsc_sp44 ^ multm_reduce_mulsc_shrsc_cp44;
  assign multm_reduce_mulsc_shrsc_sq45 = multm_reduce_mulsc_shrsc_sp45 ^ multm_reduce_mulsc_shrsc_cp45;
  assign multm_reduce_mulsc_shrsc_sq46 = multm_reduce_mulsc_shrsc_sp46 ^ multm_reduce_mulsc_shrsc_cp46;
  assign multm_reduce_mulsc_shrsc_sq47 = multm_reduce_mulsc_shrsc_sp47 ^ multm_reduce_mulsc_shrsc_cp47;
  assign multm_reduce_mulsc_shrsc_sq48 = multm_reduce_mulsc_shrsc_sp48 ^ multm_reduce_mulsc_shrsc_cp48;
  assign multm_reduce_mulsc_shrsc_sq49 = multm_reduce_mulsc_shrsc_sp49 ^ multm_reduce_mulsc_shrsc_cp49;
  assign multm_reduce_mulsc_shrsc_sq50 = multm_reduce_mulsc_shrsc_sp50 ^ multm_reduce_mulsc_shrsc_cp50;
  assign multm_reduce_mulsc_shrsc_sq51 = multm_reduce_mulsc_shrsc_sp51 ^ multm_reduce_mulsc_shrsc_cp51;
  assign multm_reduce_mulsc_shrsc_sq52 = multm_reduce_mulsc_shrsc_sp52 ^ multm_reduce_mulsc_shrsc_cp52;
  assign multm_reduce_mulsc_shrsc_sq53 = multm_reduce_mulsc_shrsc_sp53 ^ multm_reduce_mulsc_shrsc_cp53;
  assign multm_reduce_mulsc_shrsc_sq54 = multm_reduce_mulsc_shrsc_sp54 ^ multm_reduce_mulsc_shrsc_cp54;
  assign multm_reduce_mulsc_shrsc_sq55 = multm_reduce_mulsc_shrsc_sp55 ^ multm_reduce_mulsc_shrsc_cp55;
  assign multm_reduce_mulsc_shrsc_sq56 = multm_reduce_mulsc_shrsc_sp56 ^ multm_reduce_mulsc_shrsc_cp56;
  assign multm_reduce_mulsc_shrsc_sq57 = multm_reduce_mulsc_shrsc_sp57 ^ multm_reduce_mulsc_shrsc_cp57;
  assign multm_reduce_mulsc_shrsc_sq58 = multm_reduce_mulsc_shrsc_sp58 ^ multm_reduce_mulsc_shrsc_cp58;
  assign multm_reduce_mulsc_shrsc_sq59 = multm_reduce_mulsc_shrsc_sp59 ^ multm_reduce_mulsc_shrsc_cp59;
  assign multm_reduce_mulsc_shrsc_sq60 = multm_reduce_mulsc_shrsc_sp60 ^ multm_reduce_mulsc_shrsc_cp60;
  assign multm_reduce_mulsc_shrsc_sq61 = multm_reduce_mulsc_shrsc_sp61 ^ multm_reduce_mulsc_shrsc_cp61;
  assign multm_reduce_mulsc_shrsc_sq62 = multm_reduce_mulsc_shrsc_sp62 ^ multm_reduce_mulsc_shrsc_cp62;
  assign multm_reduce_mulsc_shrsc_sq63 = multm_reduce_mulsc_shrsc_sp63 ^ multm_reduce_mulsc_shrsc_cp63;
  assign multm_reduce_mulsc_shrsc_sq64 = multm_reduce_mulsc_shrsc_sp64 ^ multm_reduce_mulsc_shrsc_cp64;
  assign multm_reduce_mulsc_shrsc_sq65 = multm_reduce_mulsc_shrsc_sp65 ^ multm_reduce_mulsc_shrsc_cp65;
  assign multm_reduce_mulsc_shrsc_sq66 = multm_reduce_mulsc_shrsc_sp66 ^ multm_reduce_mulsc_shrsc_cp66;
  assign multm_reduce_mulsc_shrsc_sq67 = multm_reduce_mulsc_shrsc_sp67 ^ multm_reduce_mulsc_shrsc_cp67;
  assign multm_reduce_mulsc_shrsc_sq68 = multm_reduce_mulsc_shrsc_sp68 ^ multm_reduce_mulsc_shrsc_cp68;
  assign multm_reduce_mulsc_shrsc_sq69 = multm_reduce_mulsc_shrsc_sp69 ^ multm_reduce_mulsc_shrsc_cp69;
  assign multm_reduce_mulsc_shrsc_sq70 = multm_reduce_mulsc_shrsc_sp70 ^ multm_reduce_mulsc_shrsc_cp70;
  assign multm_reduce_mulsc_shrsc_sq71 = multm_reduce_mulsc_shrsc_sp71 ^ multm_reduce_mulsc_shrsc_cp71;
  assign multm_reduce_mulsc_shrsc_sq72 = multm_reduce_mulsc_shrsc_sp72 ^ multm_reduce_mulsc_shrsc_cp72;
  assign multm_reduce_mulsc_shrsc_sq73 = multm_reduce_mulsc_shrsc_sp73 ^ multm_reduce_mulsc_shrsc_cp73;
  assign multm_reduce_mulsc_shrsc_sq74 = multm_reduce_mulsc_shrsc_sp74 ^ multm_reduce_mulsc_shrsc_cp74;
  assign multm_reduce_mulsc_shrsc_sq75 = multm_reduce_mulsc_shrsc_sp75 ^ multm_reduce_mulsc_shrsc_cp75;
  assign multm_reduce_mulsc_shrsc_sq76 = multm_reduce_mulsc_shrsc_sp76 ^ multm_reduce_mulsc_shrsc_cp76;
  assign multm_reduce_mulsc_shrsc_sq77 = multm_reduce_mulsc_shrsc_sp77 ^ multm_reduce_mulsc_shrsc_cp77;
  assign multm_reduce_mulsc_shrsc_sq78 = multm_reduce_mulsc_shrsc_sp78 ^ multm_reduce_mulsc_shrsc_cp78;
  assign multm_reduce_mulsc_shrsc_sq79 = multm_reduce_mulsc_shrsc_sp79 ^ multm_reduce_mulsc_shrsc_cp79;
  assign multm_reduce_mulsc_shrsc_sq80 = multm_reduce_mulsc_shrsc_sp80 ^ multm_reduce_mulsc_shrsc_cp80;
  assign multm_reduce_mulsc_shrsc_sq81 = multm_reduce_mulsc_shrsc_sp81 ^ multm_reduce_mulsc_shrsc_cp81;
  assign multm_reduce_mulsc_shrsc_sq82 = multm_reduce_mulsc_shrsc_sp82 ^ multm_reduce_mulsc_shrsc_cp82;
  assign multm_reduce_mulsc_shrsc_sq83 = multm_reduce_mulsc_shrsc_sp83 ^ multm_reduce_mulsc_shrsc_cp83;
  assign multm_reduce_mulsc_shrsc_sq84 = multm_reduce_mulsc_shrsc_sp84 ^ multm_reduce_mulsc_shrsc_cp84;
  assign multm_reduce_mulsc_shrsc_sq85 = multm_reduce_mulsc_shrsc_sp85 ^ multm_reduce_mulsc_shrsc_cp85;
  assign multm_reduce_mulsc_shrsc_sq86 = multm_reduce_mulsc_shrsc_sp86 ^ multm_reduce_mulsc_shrsc_cp86;
  assign multm_reduce_mulsc_shrsc_sq87 = multm_reduce_mulsc_shrsc_sp87 ^ multm_reduce_mulsc_shrsc_cp87;
  assign multm_reduce_mulsc_shrsc_sq88 = multm_reduce_mulsc_shrsc_sp88 ^ multm_reduce_mulsc_shrsc_cp88;
  assign multm_reduce_mulsc_shrsc_sq89 = multm_reduce_mulsc_shrsc_sp89 ^ multm_reduce_mulsc_shrsc_cp89;
  assign multm_reduce_mulsc_shrsc_sq90 = multm_reduce_mulsc_shrsc_sp90 ^ multm_reduce_mulsc_shrsc_cp90;
  assign multm_reduce_mulsc_shrsc_sq91 = multm_reduce_mulsc_shrsc_sp91 ^ multm_reduce_mulsc_shrsc_cp91;
  assign multm_reduce_mulsc_shrsc_sq92 = multm_reduce_mulsc_shrsc_sp92 ^ multm_reduce_mulsc_shrsc_cp92;
  assign multm_reduce_mulsc_shrsc_sq93 = multm_reduce_mulsc_shrsc_sp93 ^ multm_reduce_mulsc_shrsc_cp93;
  assign multm_reduce_mulsc_shrsc_sq94 = multm_reduce_mulsc_shrsc_sp94 ^ multm_reduce_mulsc_shrsc_cp94;
  assign multm_reduce_mulsc_shrsc_sq95 = multm_reduce_mulsc_shrsc_sp95 ^ multm_reduce_mulsc_shrsc_cp95;
  assign multm_reduce_mulsc_shrsc_sq96 = multm_reduce_mulsc_shrsc_sp96 ^ multm_reduce_mulsc_shrsc_cp96;
  assign multm_reduce_mulsc_shrsc_sq97 = multm_reduce_mulsc_shrsc_sp97 ^ multm_reduce_mulsc_shrsc_cp97;
  assign multm_reduce_mulsc_shrsc_sq98 = multm_reduce_mulsc_shrsc_sp98 ^ multm_reduce_mulsc_shrsc_cp98;
  assign multm_reduce_mulsc_shrsc_sq99 = multm_reduce_mulsc_shrsc_sp99 ^ multm_reduce_mulsc_shrsc_cp99;
  assign multm_reduce_mulsc_shrsc_sq100 = multm_reduce_mulsc_shrsc_sp100 ^ multm_reduce_mulsc_shrsc_cp100;
  assign multm_reduce_mulsc_shrsc_sq101 = multm_reduce_mulsc_shrsc_sp101 ^ multm_reduce_mulsc_shrsc_cp101;
  assign multm_reduce_mulsc_shrsc_sq102 = multm_reduce_mulsc_shrsc_sp102 ^ multm_reduce_mulsc_shrsc_cp102;
  assign multm_reduce_mulsc_shrsc_sq103 = multm_reduce_mulsc_shrsc_sp103 ^ multm_reduce_mulsc_shrsc_cp103;
  assign multm_reduce_mulsc_shrsc_sq104 = multm_reduce_mulsc_shrsc_sp104 ^ multm_reduce_mulsc_shrsc_cp104;
  assign multm_reduce_mulsc_shrsc_sq105 = multm_reduce_mulsc_shrsc_sp105 ^ multm_reduce_mulsc_shrsc_cp105;
  assign multm_reduce_mulsc_shrsc_sq106 = multm_reduce_mulsc_shrsc_sp106 ^ multm_reduce_mulsc_shrsc_cp106;
  assign multm_reduce_mulsc_shrsc_sq107 = multm_reduce_mulsc_shrsc_sp107 ^ multm_reduce_mulsc_shrsc_cp107;
  assign multm_reduce_mulsc_shrsc_sq108 = multm_reduce_mulsc_shrsc_sp108 ^ multm_reduce_mulsc_shrsc_cp108;
  assign multm_reduce_mulsc_shrsc_sq109 = multm_reduce_mulsc_shrsc_sp109 ^ multm_reduce_mulsc_shrsc_cp109;
  assign multm_reduce_mulsc_shrsc_sq110 = multm_reduce_mulsc_shrsc_sp110 ^ multm_reduce_mulsc_shrsc_cp110;
  assign multm_reduce_mulsc_shrsc_sq111 = multm_reduce_mulsc_shrsc_sp111 ^ multm_reduce_mulsc_shrsc_cp111;
  assign multm_reduce_mulsc_shrsc_sq112 = multm_reduce_mulsc_shrsc_sp112 ^ multm_reduce_mulsc_shrsc_cp112;
  assign multm_reduce_mulsc_shrsc_sq113 = multm_reduce_mulsc_shrsc_sp113 ^ multm_reduce_mulsc_shrsc_cp113;
  assign multm_reduce_mulsc_shrsc_sq114 = multm_reduce_mulsc_shrsc_sp114 ^ multm_reduce_mulsc_shrsc_cp114;
  assign multm_reduce_mulsc_shrsc_sq115 = multm_reduce_mulsc_shrsc_sp115 ^ multm_reduce_mulsc_shrsc_cp115;
  assign multm_reduce_mulsc_shrsc_sq116 = multm_reduce_mulsc_shrsc_sp116 ^ multm_reduce_mulsc_shrsc_cp116;
  assign multm_reduce_mulsc_shrsc_sq117 = multm_reduce_mulsc_shrsc_sp117 ^ multm_reduce_mulsc_shrsc_cp117;
  assign multm_reduce_mulsc_shrsc_sq118 = multm_reduce_mulsc_shrsc_sp118 ^ multm_reduce_mulsc_shrsc_cp118;
  assign multm_reduce_mulsc_shrsc_sq119 = multm_reduce_mulsc_shrsc_sp119 ^ multm_reduce_mulsc_shrsc_cp119;
  assign multm_reduce_mulsc_shrsc_sq120 = multm_reduce_mulsc_shrsc_sp120 ^ multm_reduce_mulsc_shrsc_cp120;
  assign multm_reduce_mulsc_shrsc_sq121 = multm_reduce_mulsc_shrsc_sp121 ^ multm_reduce_mulsc_shrsc_cp121;
  assign multm_reduce_mulsc_shrsc_sq122 = multm_reduce_mulsc_shrsc_sp122 ^ multm_reduce_mulsc_shrsc_cp122;
  assign multm_reduce_mulsc_shrsc_sq123 = multm_reduce_mulsc_shrsc_sp123 ^ multm_reduce_mulsc_shrsc_cp123;
  assign multm_reduce_mulsc_shrsc_sq124 = multm_reduce_mulsc_shrsc_sp124 ^ multm_reduce_mulsc_shrsc_cp124;
  assign multm_reduce_mulsc_shrsc_sq125 = multm_reduce_mulsc_shrsc_sp125 ^ multm_reduce_mulsc_shrsc_cp125;
  assign multm_reduce_mulsc_shrsc_sq126 = multm_reduce_mulsc_shrsc_sp126 ^ multm_reduce_mulsc_shrsc_cp126;
  assign multm_reduce_mulsc_shrsc_sq127 = multm_reduce_mulsc_shrsc_sp127 ^ multm_reduce_mulsc_shrsc_cp127;
  assign multm_reduce_mulsc_shrsc_sq128 = multm_reduce_mulsc_shrsc_sp128 ^ multm_reduce_mulsc_shrsc_cp128;
  assign multm_reduce_mulsc_shrsc_sq129 = multm_reduce_mulsc_shrsc_sp129 ^ multm_reduce_mulsc_shrsc_cp129;
  assign multm_reduce_mulsc_shrsc_sq130 = multm_reduce_mulsc_shrsc_sp130 ^ multm_reduce_mulsc_shrsc_cp130;
  assign multm_reduce_mulsc_shrsc_sq131 = multm_reduce_mulsc_shrsc_sp131 ^ multm_reduce_mulsc_shrsc_cp131;
  assign multm_reduce_mulsc_shrsc_sq132 = multm_reduce_mulsc_shrsc_sp132 ^ multm_reduce_mulsc_shrsc_cp132;
  assign multm_reduce_mulsc_shrsc_sq133 = multm_reduce_mulsc_shrsc_sp133 ^ multm_reduce_mulsc_shrsc_cp133;
  assign multm_reduce_mulsc_shrsc_sq134 = multm_reduce_mulsc_shrsc_sp134 ^ multm_reduce_mulsc_shrsc_cp134;
  assign multm_reduce_mulsc_shrsc_sq135 = multm_reduce_mulsc_shrsc_sp135 ^ multm_reduce_mulsc_shrsc_cp135;
  assign multm_reduce_mulsc_shrsc_sq136 = multm_reduce_mulsc_shrsc_sp136 ^ multm_reduce_mulsc_shrsc_cp136;
  assign multm_reduce_mulsc_shrsc_sq137 = multm_reduce_mulsc_shrsc_sp137 ^ multm_reduce_mulsc_shrsc_cp137;
  assign multm_reduce_mulsc_shrsc_sq138 = multm_reduce_mulsc_shrsc_sp138 ^ multm_reduce_mulsc_shrsc_cp138;
  assign multm_reduce_mulsc_shrsc_sq139 = multm_reduce_mulsc_shrsc_sp139 ^ multm_reduce_mulsc_shrsc_cp139;
  assign multm_reduce_mulsc_shrsc_sq140 = multm_reduce_mulsc_shrsc_sp140 ^ multm_reduce_mulsc_shrsc_cp140;
  assign multm_reduce_mulsc_shrsc_sq141 = multm_reduce_mulsc_shrsc_sp141 ^ multm_reduce_mulsc_shrsc_cp141;
  assign multm_reduce_mulsc_shrsc_sq142 = multm_reduce_mulsc_shrsc_sp142 ^ multm_reduce_mulsc_shrsc_cp142;
  assign multm_reduce_mulsc_shrsc_sq143 = multm_reduce_mulsc_shrsc_sp143 ^ multm_reduce_mulsc_shrsc_cp143;
  assign multm_reduce_mulsc_shrsc_sq144 = multm_reduce_mulsc_shrsc_sp144 ^ multm_reduce_mulsc_shrsc_cp144;
  assign multm_reduce_mulsc_shrsc_sq145 = multm_reduce_mulsc_shrsc_sp145 ^ multm_reduce_mulsc_shrsc_cp145;
  assign multm_reduce_mulsc_shrsc_sq146 = multm_reduce_mulsc_shrsc_sp146 ^ multm_reduce_mulsc_shrsc_cp146;
  assign multm_reduce_mulsc_shrsc_sq147 = multm_reduce_mulsc_shrsc_sp147 ^ multm_reduce_mulsc_shrsc_cp147;
  assign multm_reduce_mulsc_shrsc_sq148 = multm_reduce_mulsc_shrsc_sp148 ^ multm_reduce_mulsc_shrsc_cp148;
  assign multm_reduce_mulsc_shrsc_sq149 = multm_reduce_mulsc_shrsc_sp149 ^ multm_reduce_mulsc_shrsc_cp149;
  assign multm_reduce_mulsc_shrsc_sq150 = multm_reduce_mulsc_shrsc_sp150 ^ multm_reduce_mulsc_shrsc_cp150;
  assign multm_reduce_mulsc_shrsc_sq151 = multm_reduce_mulsc_shrsc_sp151 ^ multm_reduce_mulsc_shrsc_cp151;
  assign multm_reduce_mulsc_shrsc_sq152 = multm_reduce_mulsc_shrsc_sp152 ^ multm_reduce_mulsc_shrsc_cp152;
  assign multm_reduce_mulsc_shrsc_sq153 = multm_reduce_mulsc_shrsc_sp153 ^ multm_reduce_mulsc_shrsc_cp153;
  assign multm_reduce_mulsc_shrsc_sq154 = multm_reduce_mulsc_shrsc_sp154 ^ multm_reduce_mulsc_shrsc_cp154;
  assign multm_reduce_mulsc_shrsc_sq155 = multm_reduce_mulsc_shrsc_sp155 ^ multm_reduce_mulsc_shrsc_cp155;
  assign multm_reduce_mulsc_shrsc_sq156 = multm_reduce_mulsc_shrsc_sp156 ^ multm_reduce_mulsc_shrsc_cp156;
  assign multm_reduce_mulsc_shrsc_sq157 = multm_reduce_mulsc_shrsc_sp157 ^ multm_reduce_mulsc_shrsc_cp157;
  assign multm_reduce_mulsc_shrsc_sq158 = multm_reduce_mulsc_shrsc_sp158 ^ multm_reduce_mulsc_shrsc_cp158;
  assign multm_reduce_mulsc_shrsc_sq159 = multm_reduce_mulsc_shrsc_sp159 ^ multm_reduce_mulsc_shrsc_cp159;
  assign multm_reduce_mulsc_shrsc_sq160 = multm_reduce_mulsc_shrsc_sp160 ^ multm_reduce_mulsc_shrsc_cp160;
  assign multm_reduce_mulsc_shrsc_sq161 = multm_reduce_mulsc_shrsc_sp161 ^ multm_reduce_mulsc_shrsc_cp161;
  assign multm_reduce_mulsc_shrsc_sq162 = multm_reduce_mulsc_shrsc_sp162 ^ multm_reduce_mulsc_shrsc_cp162;
  assign multm_reduce_mulsc_shrsc_sq163 = multm_reduce_mulsc_shrsc_sp163 ^ multm_reduce_mulsc_shrsc_cp163;
  assign multm_reduce_mulsc_shrsc_sq164 = multm_reduce_mulsc_shrsc_sp164 ^ multm_reduce_mulsc_shrsc_cp164;
  assign multm_reduce_mulsc_shrsc_sq165 = multm_reduce_mulsc_shrsc_sp165 ^ multm_reduce_mulsc_shrsc_cp165;
  assign multm_reduce_mulsc_shrsc_sq166 = multm_reduce_mulsc_shrsc_sp166 ^ multm_reduce_mulsc_shrsc_cp166;
  assign multm_reduce_mulsc_shrsc_sq167 = multm_reduce_mulsc_shrsc_sp167 ^ multm_reduce_mulsc_shrsc_cp167;
  assign multm_reduce_mulsc_shrsc_sq168 = multm_reduce_mulsc_shrsc_sp168 ^ multm_reduce_mulsc_shrsc_cp168;
  assign multm_reduce_mulsc_shrsc_sq169 = multm_reduce_mulsc_shrsc_sp169 ^ multm_reduce_mulsc_shrsc_cp169;
  assign multm_reduce_mulsc_shrsc_sq170 = multm_reduce_mulsc_shrsc_sp170 ^ multm_reduce_mulsc_shrsc_cp170;
  assign multm_reduce_mulsc_shrsc_sq171 = multm_reduce_mulsc_shrsc_sp171 ^ multm_reduce_mulsc_shrsc_cp171;
  assign multm_reduce_mulsc_shrsc_sq172 = multm_reduce_mulsc_shrsc_sp172 ^ multm_reduce_mulsc_shrsc_cp172;
  assign multm_reduce_mulsc_shrsc_sq173 = multm_reduce_mulsc_shrsc_sp173 ^ multm_reduce_mulsc_shrsc_cp173;
  assign multm_reduce_mulsc_shrsc_sq174 = multm_reduce_mulsc_shrsc_sp174 ^ multm_reduce_mulsc_shrsc_cp174;
  assign multm_reduce_mulsc_shrsc_sq175 = multm_reduce_mulsc_shrsc_sp175 ^ multm_reduce_mulsc_shrsc_cp175;
  assign multm_reduce_mulsc_shrsc_sq176 = multm_reduce_mulsc_shrsc_sp176 ^ multm_reduce_mulsc_shrsc_cp176;
  assign multm_reduce_mulsc_shrsc_sq177 = multm_reduce_mulsc_shrsc_sp177 ^ multm_reduce_mulsc_shrsc_cp177;
  assign multm_reduce_mulsc_shrsc_sq178 = multm_reduce_mulsc_shrsc_sp178 ^ multm_reduce_mulsc_shrsc_cp178;
  assign multm_reduce_mulsc_shrsc_sq179 = multm_reduce_mulsc_shrsc_sp179 ^ multm_reduce_mulsc_shrsc_cp179;
  assign multm_reduce_mulsc_shrsc_sq180 = multm_reduce_mulsc_shrsc_sp180 ^ multm_reduce_mulsc_shrsc_cp180;
  assign multm_reduce_mulsc_shrsc_sq181 = multm_reduce_mulsc_shrsc_sp181 ^ multm_reduce_mulsc_shrsc_cp181;
  assign multm_reduce_mulsc_shrsc_sq182 = multm_reduce_mulsc_shrsc_sp182 ^ multm_reduce_mulsc_shrsc_cp182;
  assign multm_reduce_mulsc_shrsc_sr0 = sadd ? ys1_o : multm_reduce_mulsc_shrsc_sq1;
  assign multm_reduce_mulsc_shrsc_sr1 = sadd ? ys2_o : multm_reduce_mulsc_shrsc_sq2;
  assign multm_reduce_mulsc_shrsc_sr2 = sadd ? ys3_o : multm_reduce_mulsc_shrsc_sq3;
  assign multm_reduce_mulsc_shrsc_sr3 = sadd ? ys4_o : multm_reduce_mulsc_shrsc_sq4;
  assign multm_reduce_mulsc_shrsc_sr4 = sadd ? ys5_o : multm_reduce_mulsc_shrsc_sq5;
  assign multm_reduce_mulsc_shrsc_sr5 = sadd ? ys6_o : multm_reduce_mulsc_shrsc_sq6;
  assign multm_reduce_mulsc_shrsc_sr6 = sadd ? ys7_o : multm_reduce_mulsc_shrsc_sq7;
  assign multm_reduce_mulsc_shrsc_sr7 = sadd ? ys8_o : multm_reduce_mulsc_shrsc_sq8;
  assign multm_reduce_mulsc_shrsc_sr8 = sadd ? ys9_o : multm_reduce_mulsc_shrsc_sq9;
  assign multm_reduce_mulsc_shrsc_sr9 = sadd ? ys10_o : multm_reduce_mulsc_shrsc_sq10;
  assign multm_reduce_mulsc_shrsc_sr10 = sadd ? ys11_o : multm_reduce_mulsc_shrsc_sq11;
  assign multm_reduce_mulsc_shrsc_sr11 = sadd ? ys12_o : multm_reduce_mulsc_shrsc_sq12;
  assign multm_reduce_mulsc_shrsc_sr12 = sadd ? ys13_o : multm_reduce_mulsc_shrsc_sq13;
  assign multm_reduce_mulsc_shrsc_sr13 = sadd ? ys14_o : multm_reduce_mulsc_shrsc_sq14;
  assign multm_reduce_mulsc_shrsc_sr14 = sadd ? ys15_o : multm_reduce_mulsc_shrsc_sq15;
  assign multm_reduce_mulsc_shrsc_sr15 = sadd ? ys16_o : multm_reduce_mulsc_shrsc_sq16;
  assign multm_reduce_mulsc_shrsc_sr16 = sadd ? ys17_o : multm_reduce_mulsc_shrsc_sq17;
  assign multm_reduce_mulsc_shrsc_sr17 = sadd ? ys18_o : multm_reduce_mulsc_shrsc_sq18;
  assign multm_reduce_mulsc_shrsc_sr18 = sadd ? ys19_o : multm_reduce_mulsc_shrsc_sq19;
  assign multm_reduce_mulsc_shrsc_sr19 = sadd ? ys20_o : multm_reduce_mulsc_shrsc_sq20;
  assign multm_reduce_mulsc_shrsc_sr20 = sadd ? ys21_o : multm_reduce_mulsc_shrsc_sq21;
  assign multm_reduce_mulsc_shrsc_sr21 = sadd ? ys22_o : multm_reduce_mulsc_shrsc_sq22;
  assign multm_reduce_mulsc_shrsc_sr22 = sadd ? ys23_o : multm_reduce_mulsc_shrsc_sq23;
  assign multm_reduce_mulsc_shrsc_sr23 = sadd ? ys24_o : multm_reduce_mulsc_shrsc_sq24;
  assign multm_reduce_mulsc_shrsc_sr24 = sadd ? ys25_o : multm_reduce_mulsc_shrsc_sq25;
  assign multm_reduce_mulsc_shrsc_sr25 = sadd ? ys26_o : multm_reduce_mulsc_shrsc_sq26;
  assign multm_reduce_mulsc_shrsc_sr26 = sadd ? ys27_o : multm_reduce_mulsc_shrsc_sq27;
  assign multm_reduce_mulsc_shrsc_sr27 = sadd ? ys28_o : multm_reduce_mulsc_shrsc_sq28;
  assign multm_reduce_mulsc_shrsc_sr28 = sadd ? ys29_o : multm_reduce_mulsc_shrsc_sq29;
  assign multm_reduce_mulsc_shrsc_sr29 = sadd ? ys30_o : multm_reduce_mulsc_shrsc_sq30;
  assign multm_reduce_mulsc_shrsc_sr30 = sadd ? ys31_o : multm_reduce_mulsc_shrsc_sq31;
  assign multm_reduce_mulsc_shrsc_sr31 = sadd ? ys32_o : multm_reduce_mulsc_shrsc_sq32;
  assign multm_reduce_mulsc_shrsc_sr32 = sadd ? ys33_o : multm_reduce_mulsc_shrsc_sq33;
  assign multm_reduce_mulsc_shrsc_sr33 = sadd ? ys34_o : multm_reduce_mulsc_shrsc_sq34;
  assign multm_reduce_mulsc_shrsc_sr34 = sadd ? ys35_o : multm_reduce_mulsc_shrsc_sq35;
  assign multm_reduce_mulsc_shrsc_sr35 = sadd ? ys36_o : multm_reduce_mulsc_shrsc_sq36;
  assign multm_reduce_mulsc_shrsc_sr36 = sadd ? ys37_o : multm_reduce_mulsc_shrsc_sq37;
  assign multm_reduce_mulsc_shrsc_sr37 = sadd ? ys38_o : multm_reduce_mulsc_shrsc_sq38;
  assign multm_reduce_mulsc_shrsc_sr38 = sadd ? ys39_o : multm_reduce_mulsc_shrsc_sq39;
  assign multm_reduce_mulsc_shrsc_sr39 = sadd ? ys40_o : multm_reduce_mulsc_shrsc_sq40;
  assign multm_reduce_mulsc_shrsc_sr40 = sadd ? ys41_o : multm_reduce_mulsc_shrsc_sq41;
  assign multm_reduce_mulsc_shrsc_sr41 = sadd ? ys42_o : multm_reduce_mulsc_shrsc_sq42;
  assign multm_reduce_mulsc_shrsc_sr42 = sadd ? ys43_o : multm_reduce_mulsc_shrsc_sq43;
  assign multm_reduce_mulsc_shrsc_sr43 = sadd ? ys44_o : multm_reduce_mulsc_shrsc_sq44;
  assign multm_reduce_mulsc_shrsc_sr44 = sadd ? ys45_o : multm_reduce_mulsc_shrsc_sq45;
  assign multm_reduce_mulsc_shrsc_sr45 = sadd ? ys46_o : multm_reduce_mulsc_shrsc_sq46;
  assign multm_reduce_mulsc_shrsc_sr46 = sadd ? ys47_o : multm_reduce_mulsc_shrsc_sq47;
  assign multm_reduce_mulsc_shrsc_sr47 = sadd ? ys48_o : multm_reduce_mulsc_shrsc_sq48;
  assign multm_reduce_mulsc_shrsc_sr48 = sadd ? ys49_o : multm_reduce_mulsc_shrsc_sq49;
  assign multm_reduce_mulsc_shrsc_sr49 = sadd ? ys50_o : multm_reduce_mulsc_shrsc_sq50;
  assign multm_reduce_mulsc_shrsc_sr50 = sadd ? ys51_o : multm_reduce_mulsc_shrsc_sq51;
  assign multm_reduce_mulsc_shrsc_sr51 = sadd ? ys52_o : multm_reduce_mulsc_shrsc_sq52;
  assign multm_reduce_mulsc_shrsc_sr52 = sadd ? ys53_o : multm_reduce_mulsc_shrsc_sq53;
  assign multm_reduce_mulsc_shrsc_sr53 = sadd ? ys54_o : multm_reduce_mulsc_shrsc_sq54;
  assign multm_reduce_mulsc_shrsc_sr54 = sadd ? ys55_o : multm_reduce_mulsc_shrsc_sq55;
  assign multm_reduce_mulsc_shrsc_sr55 = sadd ? ys56_o : multm_reduce_mulsc_shrsc_sq56;
  assign multm_reduce_mulsc_shrsc_sr56 = sadd ? ys57_o : multm_reduce_mulsc_shrsc_sq57;
  assign multm_reduce_mulsc_shrsc_sr57 = sadd ? ys58_o : multm_reduce_mulsc_shrsc_sq58;
  assign multm_reduce_mulsc_shrsc_sr58 = sadd ? ys59_o : multm_reduce_mulsc_shrsc_sq59;
  assign multm_reduce_mulsc_shrsc_sr59 = sadd ? ys60_o : multm_reduce_mulsc_shrsc_sq60;
  assign multm_reduce_mulsc_shrsc_sr60 = sadd ? ys61_o : multm_reduce_mulsc_shrsc_sq61;
  assign multm_reduce_mulsc_shrsc_sr61 = sadd ? ys62_o : multm_reduce_mulsc_shrsc_sq62;
  assign multm_reduce_mulsc_shrsc_sr62 = sadd ? ys63_o : multm_reduce_mulsc_shrsc_sq63;
  assign multm_reduce_mulsc_shrsc_sr63 = sadd ? ys64_o : multm_reduce_mulsc_shrsc_sq64;
  assign multm_reduce_mulsc_shrsc_sr64 = sadd ? ys65_o : multm_reduce_mulsc_shrsc_sq65;
  assign multm_reduce_mulsc_shrsc_sr65 = sadd ? ys66_o : multm_reduce_mulsc_shrsc_sq66;
  assign multm_reduce_mulsc_shrsc_sr66 = sadd ? ys67_o : multm_reduce_mulsc_shrsc_sq67;
  assign multm_reduce_mulsc_shrsc_sr67 = sadd ? ys68_o : multm_reduce_mulsc_shrsc_sq68;
  assign multm_reduce_mulsc_shrsc_sr68 = sadd ? ys69_o : multm_reduce_mulsc_shrsc_sq69;
  assign multm_reduce_mulsc_shrsc_sr69 = sadd ? ys70_o : multm_reduce_mulsc_shrsc_sq70;
  assign multm_reduce_mulsc_shrsc_sr70 = sadd ? ys71_o : multm_reduce_mulsc_shrsc_sq71;
  assign multm_reduce_mulsc_shrsc_sr71 = sadd ? ys72_o : multm_reduce_mulsc_shrsc_sq72;
  assign multm_reduce_mulsc_shrsc_sr72 = sadd ? ys73_o : multm_reduce_mulsc_shrsc_sq73;
  assign multm_reduce_mulsc_shrsc_sr73 = sadd ? ys74_o : multm_reduce_mulsc_shrsc_sq74;
  assign multm_reduce_mulsc_shrsc_sr74 = sadd ? ys75_o : multm_reduce_mulsc_shrsc_sq75;
  assign multm_reduce_mulsc_shrsc_sr75 = sadd ? ys76_o : multm_reduce_mulsc_shrsc_sq76;
  assign multm_reduce_mulsc_shrsc_sr76 = sadd ? ys77_o : multm_reduce_mulsc_shrsc_sq77;
  assign multm_reduce_mulsc_shrsc_sr77 = sadd ? ys78_o : multm_reduce_mulsc_shrsc_sq78;
  assign multm_reduce_mulsc_shrsc_sr78 = sadd ? ys79_o : multm_reduce_mulsc_shrsc_sq79;
  assign multm_reduce_mulsc_shrsc_sr79 = sadd ? ys80_o : multm_reduce_mulsc_shrsc_sq80;
  assign multm_reduce_mulsc_shrsc_sr80 = sadd ? ys81_o : multm_reduce_mulsc_shrsc_sq81;
  assign multm_reduce_mulsc_shrsc_sr81 = sadd ? ys82_o : multm_reduce_mulsc_shrsc_sq82;
  assign multm_reduce_mulsc_shrsc_sr82 = sadd ? ys83_o : multm_reduce_mulsc_shrsc_sq83;
  assign multm_reduce_mulsc_shrsc_sr83 = sadd ? ys84_o : multm_reduce_mulsc_shrsc_sq84;
  assign multm_reduce_mulsc_shrsc_sr84 = sadd ? ys85_o : multm_reduce_mulsc_shrsc_sq85;
  assign multm_reduce_mulsc_shrsc_sr85 = sadd ? ys86_o : multm_reduce_mulsc_shrsc_sq86;
  assign multm_reduce_mulsc_shrsc_sr86 = sadd ? ys87_o : multm_reduce_mulsc_shrsc_sq87;
  assign multm_reduce_mulsc_shrsc_sr87 = sadd ? ys88_o : multm_reduce_mulsc_shrsc_sq88;
  assign multm_reduce_mulsc_shrsc_sr88 = sadd ? ys89_o : multm_reduce_mulsc_shrsc_sq89;
  assign multm_reduce_mulsc_shrsc_sr89 = sadd ? ys90_o : multm_reduce_mulsc_shrsc_sq90;
  assign multm_reduce_mulsc_shrsc_sr90 = sadd ? ys91_o : multm_reduce_mulsc_shrsc_sq91;
  assign multm_reduce_mulsc_shrsc_sr91 = sadd ? ys92_o : multm_reduce_mulsc_shrsc_sq92;
  assign multm_reduce_mulsc_shrsc_sr92 = sadd ? ys93_o : multm_reduce_mulsc_shrsc_sq93;
  assign multm_reduce_mulsc_shrsc_sr93 = sadd ? ys94_o : multm_reduce_mulsc_shrsc_sq94;
  assign multm_reduce_mulsc_shrsc_sr94 = sadd ? ys95_o : multm_reduce_mulsc_shrsc_sq95;
  assign multm_reduce_mulsc_shrsc_sr95 = sadd ? ys96_o : multm_reduce_mulsc_shrsc_sq96;
  assign multm_reduce_mulsc_shrsc_sr96 = sadd ? ys97_o : multm_reduce_mulsc_shrsc_sq97;
  assign multm_reduce_mulsc_shrsc_sr97 = sadd ? ys98_o : multm_reduce_mulsc_shrsc_sq98;
  assign multm_reduce_mulsc_shrsc_sr98 = sadd ? ys99_o : multm_reduce_mulsc_shrsc_sq99;
  assign multm_reduce_mulsc_shrsc_sr99 = sadd ? ys100_o : multm_reduce_mulsc_shrsc_sq100;
  assign multm_reduce_mulsc_shrsc_sr100 = sadd ? ys101_o : multm_reduce_mulsc_shrsc_sq101;
  assign multm_reduce_mulsc_shrsc_sr101 = sadd ? ys102_o : multm_reduce_mulsc_shrsc_sq102;
  assign multm_reduce_mulsc_shrsc_sr102 = sadd ? ys103_o : multm_reduce_mulsc_shrsc_sq103;
  assign multm_reduce_mulsc_shrsc_sr103 = sadd ? ys104_o : multm_reduce_mulsc_shrsc_sq104;
  assign multm_reduce_mulsc_shrsc_sr104 = sadd ? ys105_o : multm_reduce_mulsc_shrsc_sq105;
  assign multm_reduce_mulsc_shrsc_sr105 = sadd ? ys106_o : multm_reduce_mulsc_shrsc_sq106;
  assign multm_reduce_mulsc_shrsc_sr106 = sadd ? ys107_o : multm_reduce_mulsc_shrsc_sq107;
  assign multm_reduce_mulsc_shrsc_sr107 = sadd ? ys108_o : multm_reduce_mulsc_shrsc_sq108;
  assign multm_reduce_mulsc_shrsc_sr108 = sadd ? ys109_o : multm_reduce_mulsc_shrsc_sq109;
  assign multm_reduce_mulsc_shrsc_sr109 = sadd ? ys110_o : multm_reduce_mulsc_shrsc_sq110;
  assign multm_reduce_mulsc_shrsc_sr110 = sadd ? ys111_o : multm_reduce_mulsc_shrsc_sq111;
  assign multm_reduce_mulsc_shrsc_sr111 = sadd ? ys112_o : multm_reduce_mulsc_shrsc_sq112;
  assign multm_reduce_mulsc_shrsc_sr112 = sadd ? ys113_o : multm_reduce_mulsc_shrsc_sq113;
  assign multm_reduce_mulsc_shrsc_sr113 = sadd ? ys114_o : multm_reduce_mulsc_shrsc_sq114;
  assign multm_reduce_mulsc_shrsc_sr114 = sadd ? ys115_o : multm_reduce_mulsc_shrsc_sq115;
  assign multm_reduce_mulsc_shrsc_sr115 = sadd ? ys116_o : multm_reduce_mulsc_shrsc_sq116;
  assign multm_reduce_mulsc_shrsc_sr116 = sadd ? ys117_o : multm_reduce_mulsc_shrsc_sq117;
  assign multm_reduce_mulsc_shrsc_sr117 = sadd ? ys118_o : multm_reduce_mulsc_shrsc_sq118;
  assign multm_reduce_mulsc_shrsc_sr118 = sadd ? ys119_o : multm_reduce_mulsc_shrsc_sq119;
  assign multm_reduce_mulsc_shrsc_sr119 = sadd ? ys120_o : multm_reduce_mulsc_shrsc_sq120;
  assign multm_reduce_mulsc_shrsc_sr120 = sadd ? ys121_o : multm_reduce_mulsc_shrsc_sq121;
  assign multm_reduce_mulsc_shrsc_sr121 = sadd ? ys122_o : multm_reduce_mulsc_shrsc_sq122;
  assign multm_reduce_mulsc_shrsc_sr122 = sadd ? ys123_o : multm_reduce_mulsc_shrsc_sq123;
  assign multm_reduce_mulsc_shrsc_sr123 = sadd ? ys124_o : multm_reduce_mulsc_shrsc_sq124;
  assign multm_reduce_mulsc_shrsc_sr124 = sadd ? ys125_o : multm_reduce_mulsc_shrsc_sq125;
  assign multm_reduce_mulsc_shrsc_sr125 = sadd ? ys126_o : multm_reduce_mulsc_shrsc_sq126;
  assign multm_reduce_mulsc_shrsc_sr126 = sadd ? ys127_o : multm_reduce_mulsc_shrsc_sq127;
  assign multm_reduce_mulsc_shrsc_sr127 = sadd ? ys128_o : multm_reduce_mulsc_shrsc_sq128;
  assign multm_reduce_mulsc_shrsc_sr128 = sadd ? ys129_o : multm_reduce_mulsc_shrsc_sq129;
  assign multm_reduce_mulsc_shrsc_sr129 = sadd ? ys130_o : multm_reduce_mulsc_shrsc_sq130;
  assign multm_reduce_mulsc_shrsc_sr130 = sadd ? ys131_o : multm_reduce_mulsc_shrsc_sq131;
  assign multm_reduce_mulsc_shrsc_sr131 = sadd ? ys132_o : multm_reduce_mulsc_shrsc_sq132;
  assign multm_reduce_mulsc_shrsc_sr132 = sadd ? ys133_o : multm_reduce_mulsc_shrsc_sq133;
  assign multm_reduce_mulsc_shrsc_sr133 = sadd ? ys134_o : multm_reduce_mulsc_shrsc_sq134;
  assign multm_reduce_mulsc_shrsc_sr134 = sadd ? ys135_o : multm_reduce_mulsc_shrsc_sq135;
  assign multm_reduce_mulsc_shrsc_sr135 = sadd ? ys136_o : multm_reduce_mulsc_shrsc_sq136;
  assign multm_reduce_mulsc_shrsc_sr136 = sadd ? ys137_o : multm_reduce_mulsc_shrsc_sq137;
  assign multm_reduce_mulsc_shrsc_sr137 = sadd ? ys138_o : multm_reduce_mulsc_shrsc_sq138;
  assign multm_reduce_mulsc_shrsc_sr138 = sadd ? ys139_o : multm_reduce_mulsc_shrsc_sq139;
  assign multm_reduce_mulsc_shrsc_sr139 = sadd ? ys140_o : multm_reduce_mulsc_shrsc_sq140;
  assign multm_reduce_mulsc_shrsc_sr140 = sadd ? ys141_o : multm_reduce_mulsc_shrsc_sq141;
  assign multm_reduce_mulsc_shrsc_sr141 = sadd ? ys142_o : multm_reduce_mulsc_shrsc_sq142;
  assign multm_reduce_mulsc_shrsc_sr142 = sadd ? ys143_o : multm_reduce_mulsc_shrsc_sq143;
  assign multm_reduce_mulsc_shrsc_sr143 = sadd ? ys144_o : multm_reduce_mulsc_shrsc_sq144;
  assign multm_reduce_mulsc_shrsc_sr144 = sadd ? ys145_o : multm_reduce_mulsc_shrsc_sq145;
  assign multm_reduce_mulsc_shrsc_sr145 = sadd ? ys146_o : multm_reduce_mulsc_shrsc_sq146;
  assign multm_reduce_mulsc_shrsc_sr146 = sadd ? ys147_o : multm_reduce_mulsc_shrsc_sq147;
  assign multm_reduce_mulsc_shrsc_sr147 = sadd ? ys148_o : multm_reduce_mulsc_shrsc_sq148;
  assign multm_reduce_mulsc_shrsc_sr148 = sadd ? ys149_o : multm_reduce_mulsc_shrsc_sq149;
  assign multm_reduce_mulsc_shrsc_sr149 = sadd ? ys150_o : multm_reduce_mulsc_shrsc_sq150;
  assign multm_reduce_mulsc_shrsc_sr150 = sadd ? ys151_o : multm_reduce_mulsc_shrsc_sq151;
  assign multm_reduce_mulsc_shrsc_sr151 = sadd ? ys152_o : multm_reduce_mulsc_shrsc_sq152;
  assign multm_reduce_mulsc_shrsc_sr152 = sadd ? ys153_o : multm_reduce_mulsc_shrsc_sq153;
  assign multm_reduce_mulsc_shrsc_sr153 = sadd ? ys154_o : multm_reduce_mulsc_shrsc_sq154;
  assign multm_reduce_mulsc_shrsc_sr154 = sadd ? ys155_o : multm_reduce_mulsc_shrsc_sq155;
  assign multm_reduce_mulsc_shrsc_sr155 = sadd ? ys156_o : multm_reduce_mulsc_shrsc_sq156;
  assign multm_reduce_mulsc_shrsc_sr156 = sadd ? ys157_o : multm_reduce_mulsc_shrsc_sq157;
  assign multm_reduce_mulsc_shrsc_sr157 = sadd ? ys158_o : multm_reduce_mulsc_shrsc_sq158;
  assign multm_reduce_mulsc_shrsc_sr158 = sadd ? ys159_o : multm_reduce_mulsc_shrsc_sq159;
  assign multm_reduce_mulsc_shrsc_sr159 = sadd ? ys160_o : multm_reduce_mulsc_shrsc_sq160;
  assign multm_reduce_mulsc_shrsc_sr160 = sadd ? ys161_o : multm_reduce_mulsc_shrsc_sq161;
  assign multm_reduce_mulsc_shrsc_sr161 = sadd ? ys162_o : multm_reduce_mulsc_shrsc_sq162;
  assign multm_reduce_mulsc_shrsc_sr162 = sadd ? ys163_o : multm_reduce_mulsc_shrsc_sq163;
  assign multm_reduce_mulsc_shrsc_sr163 = sadd ? ys164_o : multm_reduce_mulsc_shrsc_sq164;
  assign multm_reduce_mulsc_shrsc_sr164 = sadd ? ys165_o : multm_reduce_mulsc_shrsc_sq165;
  assign multm_reduce_mulsc_shrsc_sr165 = sadd ? ys166_o : multm_reduce_mulsc_shrsc_sq166;
  assign multm_reduce_mulsc_shrsc_sr166 = sadd ? ys167_o : multm_reduce_mulsc_shrsc_sq167;
  assign multm_reduce_mulsc_shrsc_sr167 = sadd ? ys168_o : multm_reduce_mulsc_shrsc_sq168;
  assign multm_reduce_mulsc_shrsc_sr168 = sadd ? ys169_o : multm_reduce_mulsc_shrsc_sq169;
  assign multm_reduce_mulsc_shrsc_sr169 = sadd ? ys170_o : multm_reduce_mulsc_shrsc_sq170;
  assign multm_reduce_mulsc_shrsc_sr170 = sadd ? ys171_o : multm_reduce_mulsc_shrsc_sq171;
  assign multm_reduce_mulsc_shrsc_sr171 = sadd ? ys172_o : multm_reduce_mulsc_shrsc_sq172;
  assign multm_reduce_mulsc_shrsc_sr172 = sadd ? ys173_o : multm_reduce_mulsc_shrsc_sq173;
  assign multm_reduce_mulsc_shrsc_sr173 = sadd ? ys174_o : multm_reduce_mulsc_shrsc_sq174;
  assign multm_reduce_mulsc_shrsc_sr174 = sadd ? ys175_o : multm_reduce_mulsc_shrsc_sq175;
  assign multm_reduce_mulsc_shrsc_sr175 = sadd ? ys176_o : multm_reduce_mulsc_shrsc_sq176;
  assign multm_reduce_mulsc_shrsc_sr176 = sadd ? ys177_o : multm_reduce_mulsc_shrsc_sq177;
  assign multm_reduce_mulsc_shrsc_sr177 = sadd ? ys178_o : multm_reduce_mulsc_shrsc_sq178;
  assign multm_reduce_mulsc_shrsc_sr178 = sadd ? ys179_o : multm_reduce_mulsc_shrsc_sq179;
  assign multm_reduce_mulsc_shrsc_sr179 = sadd ? ys180_o : multm_reduce_mulsc_shrsc_sq180;
  assign multm_reduce_mulsc_shrsc_sr180 = sadd ? ys181_o : multm_reduce_mulsc_shrsc_sq181;
  assign multm_reduce_mulsc_shrsc_sr181 = sadd ? ys182_o : multm_reduce_mulsc_shrsc_sq182;
  assign multm_reduce_mulsc_shrsc_sr182 = sadd ? ys183_o : multm_reduce_mulsc_shrsc_cp183;
  assign multm_reduce_mulsc_xb = sadd ? ys0_o : multm_reduce_mulsc_shrsc_sq0;
  assign multm_reduce_mw = multm_reduce_add3_maj3_or3_wx | multm_reduce_add3_maj3_xy;
  assign multm_reduce_or3_wx = multm_reduce_sb174 | multm_reduce_sa185;
  assign multm_reduce_pb = multm_reduce_mulsc_mulb_sq0 ^ multm_reduce_mulsc_mulb_yos0;
  assign multm_reduce_pc0 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx0 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy0;
  assign multm_reduce_pc1 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx1 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy1;
  assign multm_reduce_pc2 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx2 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy2;
  assign multm_reduce_pc3 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx3 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy3;
  assign multm_reduce_pc4 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx4 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy4;
  assign multm_reduce_pc5 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx5 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy5;
  assign multm_reduce_pc6 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx6 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy6;
  assign multm_reduce_pc7 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx7 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy7;
  assign multm_reduce_pc8 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx8 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy8;
  assign multm_reduce_pc9 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx9 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy9;
  assign multm_reduce_pc10 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx10 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy10;
  assign multm_reduce_pc11 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx11 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy11;
  assign multm_reduce_pc12 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx12 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy12;
  assign multm_reduce_pc13 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx13 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy13;
  assign multm_reduce_pc14 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx14 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy14;
  assign multm_reduce_pc15 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx15 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy15;
  assign multm_reduce_pc16 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx16 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy16;
  assign multm_reduce_pc17 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx17 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy17;
  assign multm_reduce_pc18 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx18 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy18;
  assign multm_reduce_pc19 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx19 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy19;
  assign multm_reduce_pc20 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx20 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy20;
  assign multm_reduce_pc21 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx21 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy21;
  assign multm_reduce_pc22 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx22 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy22;
  assign multm_reduce_pc23 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx23 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy23;
  assign multm_reduce_pc24 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx24 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy24;
  assign multm_reduce_pc25 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx25 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy25;
  assign multm_reduce_pc26 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx26 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy26;
  assign multm_reduce_pc27 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx27 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy27;
  assign multm_reduce_pc28 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx28 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy28;
  assign multm_reduce_pc29 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx29 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy29;
  assign multm_reduce_pc30 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx30 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy30;
  assign multm_reduce_pc31 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx31 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy31;
  assign multm_reduce_pc32 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx32 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy32;
  assign multm_reduce_pc33 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx33 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy33;
  assign multm_reduce_pc34 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx34 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy34;
  assign multm_reduce_pc35 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx35 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy35;
  assign multm_reduce_pc36 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx36 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy36;
  assign multm_reduce_pc37 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx37 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy37;
  assign multm_reduce_pc38 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx38 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy38;
  assign multm_reduce_pc39 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx39 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy39;
  assign multm_reduce_pc40 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx40 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy40;
  assign multm_reduce_pc41 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx41 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy41;
  assign multm_reduce_pc42 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx42 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy42;
  assign multm_reduce_pc43 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx43 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy43;
  assign multm_reduce_pc44 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx44 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy44;
  assign multm_reduce_pc45 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx45 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy45;
  assign multm_reduce_pc46 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx46 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy46;
  assign multm_reduce_pc47 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx47 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy47;
  assign multm_reduce_pc48 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx48 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy48;
  assign multm_reduce_pc49 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx49 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy49;
  assign multm_reduce_pc50 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx50 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy50;
  assign multm_reduce_pc51 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx51 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy51;
  assign multm_reduce_pc52 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx52 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy52;
  assign multm_reduce_pc53 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx53 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy53;
  assign multm_reduce_pc54 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx54 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy54;
  assign multm_reduce_pc55 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx55 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy55;
  assign multm_reduce_pc56 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx56 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy56;
  assign multm_reduce_pc57 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx57 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy57;
  assign multm_reduce_pc58 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx58 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy58;
  assign multm_reduce_pc59 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx59 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy59;
  assign multm_reduce_pc60 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx60 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy60;
  assign multm_reduce_pc61 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx61 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy61;
  assign multm_reduce_pc62 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx62 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy62;
  assign multm_reduce_pc63 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx63 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy63;
  assign multm_reduce_pc64 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx64 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy64;
  assign multm_reduce_pc65 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx65 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy65;
  assign multm_reduce_pc66 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx66 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy66;
  assign multm_reduce_pc67 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx67 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy67;
  assign multm_reduce_pc68 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx68 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy68;
  assign multm_reduce_pc69 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx69 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy69;
  assign multm_reduce_pc70 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx70 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy70;
  assign multm_reduce_pc71 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx71 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy71;
  assign multm_reduce_pc72 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx72 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy72;
  assign multm_reduce_pc73 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx73 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy73;
  assign multm_reduce_pc74 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx74 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy74;
  assign multm_reduce_pc75 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx75 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy75;
  assign multm_reduce_pc76 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx76 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy76;
  assign multm_reduce_pc77 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx77 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy77;
  assign multm_reduce_pc78 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx78 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy78;
  assign multm_reduce_pc79 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx79 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy79;
  assign multm_reduce_pc80 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx80 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy80;
  assign multm_reduce_pc81 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx81 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy81;
  assign multm_reduce_pc82 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx82 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy82;
  assign multm_reduce_pc83 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx83 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy83;
  assign multm_reduce_pc84 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx84 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy84;
  assign multm_reduce_pc85 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx85 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy85;
  assign multm_reduce_pc86 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx86 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy86;
  assign multm_reduce_pc87 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx87 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy87;
  assign multm_reduce_pc88 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx88 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy88;
  assign multm_reduce_pc89 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx89 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy89;
  assign multm_reduce_pc90 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx90 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy90;
  assign multm_reduce_pc91 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx91 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy91;
  assign multm_reduce_pc92 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx92 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy92;
  assign multm_reduce_pc93 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx93 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy93;
  assign multm_reduce_pc94 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx94 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy94;
  assign multm_reduce_pc95 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx95 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy95;
  assign multm_reduce_pc96 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx96 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy96;
  assign multm_reduce_pc97 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx97 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy97;
  assign multm_reduce_pc98 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx98 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy98;
  assign multm_reduce_pc99 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx99 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy99;
  assign multm_reduce_pc100 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx100 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy100;
  assign multm_reduce_pc101 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx101 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy101;
  assign multm_reduce_pc102 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx102 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy102;
  assign multm_reduce_pc103 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx103 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy103;
  assign multm_reduce_pc104 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx104 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy104;
  assign multm_reduce_pc105 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx105 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy105;
  assign multm_reduce_pc106 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx106 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy106;
  assign multm_reduce_pc107 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx107 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy107;
  assign multm_reduce_pc108 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx108 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy108;
  assign multm_reduce_pc109 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx109 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy109;
  assign multm_reduce_pc110 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx110 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy110;
  assign multm_reduce_pc111 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx111 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy111;
  assign multm_reduce_pc112 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx112 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy112;
  assign multm_reduce_pc113 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx113 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy113;
  assign multm_reduce_pc114 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx114 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy114;
  assign multm_reduce_pc115 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx115 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy115;
  assign multm_reduce_pc116 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx116 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy116;
  assign multm_reduce_pc117 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx117 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy117;
  assign multm_reduce_pc118 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx118 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy118;
  assign multm_reduce_pc119 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx119 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy119;
  assign multm_reduce_pc120 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx120 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy120;
  assign multm_reduce_pc121 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx121 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy121;
  assign multm_reduce_pc122 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx122 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy122;
  assign multm_reduce_pc123 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx123 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy123;
  assign multm_reduce_pc124 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx124 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy124;
  assign multm_reduce_pc125 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx125 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy125;
  assign multm_reduce_pc126 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx126 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy126;
  assign multm_reduce_pc127 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx127 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy127;
  assign multm_reduce_pc128 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx128 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy128;
  assign multm_reduce_pc129 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx129 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy129;
  assign multm_reduce_pc130 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx130 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy130;
  assign multm_reduce_pc131 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx131 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy131;
  assign multm_reduce_pc132 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx132 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy132;
  assign multm_reduce_pc133 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx133 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy133;
  assign multm_reduce_pc134 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx134 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy134;
  assign multm_reduce_pc135 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx135 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy135;
  assign multm_reduce_pc136 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx136 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy136;
  assign multm_reduce_pc137 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx137 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy137;
  assign multm_reduce_pc138 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx138 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy138;
  assign multm_reduce_pc139 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx139 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy139;
  assign multm_reduce_pc140 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx140 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy140;
  assign multm_reduce_pc141 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx141 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy141;
  assign multm_reduce_pc142 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx142 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy142;
  assign multm_reduce_pc143 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx143 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy143;
  assign multm_reduce_pc144 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx144 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy144;
  assign multm_reduce_pc145 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx145 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy145;
  assign multm_reduce_pc146 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx146 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy146;
  assign multm_reduce_pc147 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx147 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy147;
  assign multm_reduce_pc148 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx148 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy148;
  assign multm_reduce_pc149 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx149 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy149;
  assign multm_reduce_pc150 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx150 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy150;
  assign multm_reduce_pc151 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx151 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy151;
  assign multm_reduce_pc152 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx152 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy152;
  assign multm_reduce_pc153 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx153 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy153;
  assign multm_reduce_pc154 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx154 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy154;
  assign multm_reduce_pc155 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx155 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy155;
  assign multm_reduce_pc156 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx156 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy156;
  assign multm_reduce_pc157 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx157 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy157;
  assign multm_reduce_pc158 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx158 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy158;
  assign multm_reduce_pc159 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx159 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy159;
  assign multm_reduce_pc160 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx160 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy160;
  assign multm_reduce_pc161 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx161 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy161;
  assign multm_reduce_pc162 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx162 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy162;
  assign multm_reduce_pc163 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx163 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy163;
  assign multm_reduce_pc164 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx164 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy164;
  assign multm_reduce_pc165 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx165 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy165;
  assign multm_reduce_pc166 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx166 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy166;
  assign multm_reduce_pc167 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx167 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy167;
  assign multm_reduce_pc168 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx168 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy168;
  assign multm_reduce_pc169 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx169 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy169;
  assign multm_reduce_pc170 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx170 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy170;
  assign multm_reduce_pc171 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx171 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy171;
  assign multm_reduce_pc172 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx172 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy172;
  assign multm_reduce_pc173 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx173 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy173;
  assign multm_reduce_pc174 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx174 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy174;
  assign multm_reduce_pc175 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx175 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy175;
  assign multm_reduce_pc176 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx176 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy176;
  assign multm_reduce_pc177 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx177 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy177;
  assign multm_reduce_pc178 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx178 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy178;
  assign multm_reduce_pc179 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx179 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy179;
  assign multm_reduce_pc180 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx180 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy180;
  assign multm_reduce_pc181 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx181 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy181;
  assign multm_reduce_pc182 = multm_reduce_mulsc_mulb_add3b1_maj3b_or3b_wx182 | multm_reduce_mulsc_mulb_add3b1_maj3b_xy182;
  assign multm_reduce_pc183 = multm_reduce_mulsc_mulb_add3_maj3_or3_wx | multm_reduce_mulsc_mulb_add3_maj3_xy;
  assign multm_reduce_ps0 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx0 ^ multm_reduce_mulsc_mulb_pc0;
  assign multm_reduce_ps1 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx1 ^ multm_reduce_mulsc_mulb_pc1;
  assign multm_reduce_ps2 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx2 ^ multm_reduce_mulsc_mulb_pc2;
  assign multm_reduce_ps3 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx3 ^ multm_reduce_mulsc_mulb_pc3;
  assign multm_reduce_ps4 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx4 ^ multm_reduce_mulsc_mulb_pc4;
  assign multm_reduce_ps5 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx5 ^ multm_reduce_mulsc_mulb_pc5;
  assign multm_reduce_ps6 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx6 ^ multm_reduce_mulsc_mulb_pc6;
  assign multm_reduce_ps7 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx7 ^ multm_reduce_mulsc_mulb_pc7;
  assign multm_reduce_ps8 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx8 ^ multm_reduce_mulsc_mulb_pc8;
  assign multm_reduce_ps9 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx9 ^ multm_reduce_mulsc_mulb_pc9;
  assign multm_reduce_ps10 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx10 ^ multm_reduce_mulsc_mulb_pc10;
  assign multm_reduce_ps11 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx11 ^ multm_reduce_mulsc_mulb_pc11;
  assign multm_reduce_ps12 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx12 ^ multm_reduce_mulsc_mulb_pc12;
  assign multm_reduce_ps13 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx13 ^ multm_reduce_mulsc_mulb_pc13;
  assign multm_reduce_ps14 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx14 ^ multm_reduce_mulsc_mulb_pc14;
  assign multm_reduce_ps15 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx15 ^ multm_reduce_mulsc_mulb_pc15;
  assign multm_reduce_ps16 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx16 ^ multm_reduce_mulsc_mulb_pc16;
  assign multm_reduce_ps17 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx17 ^ multm_reduce_mulsc_mulb_pc17;
  assign multm_reduce_ps18 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx18 ^ multm_reduce_mulsc_mulb_pc18;
  assign multm_reduce_ps19 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx19 ^ multm_reduce_mulsc_mulb_pc19;
  assign multm_reduce_ps20 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx20 ^ multm_reduce_mulsc_mulb_pc20;
  assign multm_reduce_ps21 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx21 ^ multm_reduce_mulsc_mulb_pc21;
  assign multm_reduce_ps22 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx22 ^ multm_reduce_mulsc_mulb_pc22;
  assign multm_reduce_ps23 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx23 ^ multm_reduce_mulsc_mulb_pc23;
  assign multm_reduce_ps24 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx24 ^ multm_reduce_mulsc_mulb_pc24;
  assign multm_reduce_ps25 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx25 ^ multm_reduce_mulsc_mulb_pc25;
  assign multm_reduce_ps26 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx26 ^ multm_reduce_mulsc_mulb_pc26;
  assign multm_reduce_ps27 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx27 ^ multm_reduce_mulsc_mulb_pc27;
  assign multm_reduce_ps28 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx28 ^ multm_reduce_mulsc_mulb_pc28;
  assign multm_reduce_ps29 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx29 ^ multm_reduce_mulsc_mulb_pc29;
  assign multm_reduce_ps30 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx30 ^ multm_reduce_mulsc_mulb_pc30;
  assign multm_reduce_ps31 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx31 ^ multm_reduce_mulsc_mulb_pc31;
  assign multm_reduce_ps32 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx32 ^ multm_reduce_mulsc_mulb_pc32;
  assign multm_reduce_ps33 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx33 ^ multm_reduce_mulsc_mulb_pc33;
  assign multm_reduce_ps34 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx34 ^ multm_reduce_mulsc_mulb_pc34;
  assign multm_reduce_ps35 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx35 ^ multm_reduce_mulsc_mulb_pc35;
  assign multm_reduce_ps36 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx36 ^ multm_reduce_mulsc_mulb_pc36;
  assign multm_reduce_ps37 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx37 ^ multm_reduce_mulsc_mulb_pc37;
  assign multm_reduce_ps38 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx38 ^ multm_reduce_mulsc_mulb_pc38;
  assign multm_reduce_ps39 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx39 ^ multm_reduce_mulsc_mulb_pc39;
  assign multm_reduce_ps40 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx40 ^ multm_reduce_mulsc_mulb_pc40;
  assign multm_reduce_ps41 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx41 ^ multm_reduce_mulsc_mulb_pc41;
  assign multm_reduce_ps42 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx42 ^ multm_reduce_mulsc_mulb_pc42;
  assign multm_reduce_ps43 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx43 ^ multm_reduce_mulsc_mulb_pc43;
  assign multm_reduce_ps44 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx44 ^ multm_reduce_mulsc_mulb_pc44;
  assign multm_reduce_ps45 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx45 ^ multm_reduce_mulsc_mulb_pc45;
  assign multm_reduce_ps46 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx46 ^ multm_reduce_mulsc_mulb_pc46;
  assign multm_reduce_ps47 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx47 ^ multm_reduce_mulsc_mulb_pc47;
  assign multm_reduce_ps48 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx48 ^ multm_reduce_mulsc_mulb_pc48;
  assign multm_reduce_ps49 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx49 ^ multm_reduce_mulsc_mulb_pc49;
  assign multm_reduce_ps50 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx50 ^ multm_reduce_mulsc_mulb_pc50;
  assign multm_reduce_ps51 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx51 ^ multm_reduce_mulsc_mulb_pc51;
  assign multm_reduce_ps52 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx52 ^ multm_reduce_mulsc_mulb_pc52;
  assign multm_reduce_ps53 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx53 ^ multm_reduce_mulsc_mulb_pc53;
  assign multm_reduce_ps54 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx54 ^ multm_reduce_mulsc_mulb_pc54;
  assign multm_reduce_ps55 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx55 ^ multm_reduce_mulsc_mulb_pc55;
  assign multm_reduce_ps56 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx56 ^ multm_reduce_mulsc_mulb_pc56;
  assign multm_reduce_ps57 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx57 ^ multm_reduce_mulsc_mulb_pc57;
  assign multm_reduce_ps58 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx58 ^ multm_reduce_mulsc_mulb_pc58;
  assign multm_reduce_ps59 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx59 ^ multm_reduce_mulsc_mulb_pc59;
  assign multm_reduce_ps60 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx60 ^ multm_reduce_mulsc_mulb_pc60;
  assign multm_reduce_ps61 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx61 ^ multm_reduce_mulsc_mulb_pc61;
  assign multm_reduce_ps62 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx62 ^ multm_reduce_mulsc_mulb_pc62;
  assign multm_reduce_ps63 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx63 ^ multm_reduce_mulsc_mulb_pc63;
  assign multm_reduce_ps64 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx64 ^ multm_reduce_mulsc_mulb_pc64;
  assign multm_reduce_ps65 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx65 ^ multm_reduce_mulsc_mulb_pc65;
  assign multm_reduce_ps66 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx66 ^ multm_reduce_mulsc_mulb_pc66;
  assign multm_reduce_ps67 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx67 ^ multm_reduce_mulsc_mulb_pc67;
  assign multm_reduce_ps68 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx68 ^ multm_reduce_mulsc_mulb_pc68;
  assign multm_reduce_ps69 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx69 ^ multm_reduce_mulsc_mulb_pc69;
  assign multm_reduce_ps70 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx70 ^ multm_reduce_mulsc_mulb_pc70;
  assign multm_reduce_ps71 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx71 ^ multm_reduce_mulsc_mulb_pc71;
  assign multm_reduce_ps72 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx72 ^ multm_reduce_mulsc_mulb_pc72;
  assign multm_reduce_ps73 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx73 ^ multm_reduce_mulsc_mulb_pc73;
  assign multm_reduce_ps74 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx74 ^ multm_reduce_mulsc_mulb_pc74;
  assign multm_reduce_ps75 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx75 ^ multm_reduce_mulsc_mulb_pc75;
  assign multm_reduce_ps76 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx76 ^ multm_reduce_mulsc_mulb_pc76;
  assign multm_reduce_ps77 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx77 ^ multm_reduce_mulsc_mulb_pc77;
  assign multm_reduce_ps78 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx78 ^ multm_reduce_mulsc_mulb_pc78;
  assign multm_reduce_ps79 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx79 ^ multm_reduce_mulsc_mulb_pc79;
  assign multm_reduce_ps80 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx80 ^ multm_reduce_mulsc_mulb_pc80;
  assign multm_reduce_ps81 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx81 ^ multm_reduce_mulsc_mulb_pc81;
  assign multm_reduce_ps82 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx82 ^ multm_reduce_mulsc_mulb_pc82;
  assign multm_reduce_ps83 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx83 ^ multm_reduce_mulsc_mulb_pc83;
  assign multm_reduce_ps84 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx84 ^ multm_reduce_mulsc_mulb_pc84;
  assign multm_reduce_ps85 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx85 ^ multm_reduce_mulsc_mulb_pc85;
  assign multm_reduce_ps86 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx86 ^ multm_reduce_mulsc_mulb_pc86;
  assign multm_reduce_ps87 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx87 ^ multm_reduce_mulsc_mulb_pc87;
  assign multm_reduce_ps88 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx88 ^ multm_reduce_mulsc_mulb_pc88;
  assign multm_reduce_ps89 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx89 ^ multm_reduce_mulsc_mulb_pc89;
  assign multm_reduce_ps90 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx90 ^ multm_reduce_mulsc_mulb_pc90;
  assign multm_reduce_ps91 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx91 ^ multm_reduce_mulsc_mulb_pc91;
  assign multm_reduce_ps92 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx92 ^ multm_reduce_mulsc_mulb_pc92;
  assign multm_reduce_ps93 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx93 ^ multm_reduce_mulsc_mulb_pc93;
  assign multm_reduce_ps94 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx94 ^ multm_reduce_mulsc_mulb_pc94;
  assign multm_reduce_ps95 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx95 ^ multm_reduce_mulsc_mulb_pc95;
  assign multm_reduce_ps96 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx96 ^ multm_reduce_mulsc_mulb_pc96;
  assign multm_reduce_ps97 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx97 ^ multm_reduce_mulsc_mulb_pc97;
  assign multm_reduce_ps98 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx98 ^ multm_reduce_mulsc_mulb_pc98;
  assign multm_reduce_ps99 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx99 ^ multm_reduce_mulsc_mulb_pc99;
  assign multm_reduce_ps100 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx100 ^ multm_reduce_mulsc_mulb_pc100;
  assign multm_reduce_ps101 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx101 ^ multm_reduce_mulsc_mulb_pc101;
  assign multm_reduce_ps102 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx102 ^ multm_reduce_mulsc_mulb_pc102;
  assign multm_reduce_ps103 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx103 ^ multm_reduce_mulsc_mulb_pc103;
  assign multm_reduce_ps104 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx104 ^ multm_reduce_mulsc_mulb_pc104;
  assign multm_reduce_ps105 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx105 ^ multm_reduce_mulsc_mulb_pc105;
  assign multm_reduce_ps106 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx106 ^ multm_reduce_mulsc_mulb_pc106;
  assign multm_reduce_ps107 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx107 ^ multm_reduce_mulsc_mulb_pc107;
  assign multm_reduce_ps108 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx108 ^ multm_reduce_mulsc_mulb_pc108;
  assign multm_reduce_ps109 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx109 ^ multm_reduce_mulsc_mulb_pc109;
  assign multm_reduce_ps110 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx110 ^ multm_reduce_mulsc_mulb_pc110;
  assign multm_reduce_ps111 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx111 ^ multm_reduce_mulsc_mulb_pc111;
  assign multm_reduce_ps112 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx112 ^ multm_reduce_mulsc_mulb_pc112;
  assign multm_reduce_ps113 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx113 ^ multm_reduce_mulsc_mulb_pc113;
  assign multm_reduce_ps114 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx114 ^ multm_reduce_mulsc_mulb_pc114;
  assign multm_reduce_ps115 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx115 ^ multm_reduce_mulsc_mulb_pc115;
  assign multm_reduce_ps116 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx116 ^ multm_reduce_mulsc_mulb_pc116;
  assign multm_reduce_ps117 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx117 ^ multm_reduce_mulsc_mulb_pc117;
  assign multm_reduce_ps118 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx118 ^ multm_reduce_mulsc_mulb_pc118;
  assign multm_reduce_ps119 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx119 ^ multm_reduce_mulsc_mulb_pc119;
  assign multm_reduce_ps120 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx120 ^ multm_reduce_mulsc_mulb_pc120;
  assign multm_reduce_ps121 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx121 ^ multm_reduce_mulsc_mulb_pc121;
  assign multm_reduce_ps122 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx122 ^ multm_reduce_mulsc_mulb_pc122;
  assign multm_reduce_ps123 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx123 ^ multm_reduce_mulsc_mulb_pc123;
  assign multm_reduce_ps124 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx124 ^ multm_reduce_mulsc_mulb_pc124;
  assign multm_reduce_ps125 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx125 ^ multm_reduce_mulsc_mulb_pc125;
  assign multm_reduce_ps126 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx126 ^ multm_reduce_mulsc_mulb_pc126;
  assign multm_reduce_ps127 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx127 ^ multm_reduce_mulsc_mulb_pc127;
  assign multm_reduce_ps128 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx128 ^ multm_reduce_mulsc_mulb_pc128;
  assign multm_reduce_ps129 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx129 ^ multm_reduce_mulsc_mulb_pc129;
  assign multm_reduce_ps130 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx130 ^ multm_reduce_mulsc_mulb_pc130;
  assign multm_reduce_ps131 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx131 ^ multm_reduce_mulsc_mulb_pc131;
  assign multm_reduce_ps132 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx132 ^ multm_reduce_mulsc_mulb_pc132;
  assign multm_reduce_ps133 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx133 ^ multm_reduce_mulsc_mulb_pc133;
  assign multm_reduce_ps134 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx134 ^ multm_reduce_mulsc_mulb_pc134;
  assign multm_reduce_ps135 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx135 ^ multm_reduce_mulsc_mulb_pc135;
  assign multm_reduce_ps136 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx136 ^ multm_reduce_mulsc_mulb_pc136;
  assign multm_reduce_ps137 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx137 ^ multm_reduce_mulsc_mulb_pc137;
  assign multm_reduce_ps138 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx138 ^ multm_reduce_mulsc_mulb_pc138;
  assign multm_reduce_ps139 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx139 ^ multm_reduce_mulsc_mulb_pc139;
  assign multm_reduce_ps140 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx140 ^ multm_reduce_mulsc_mulb_pc140;
  assign multm_reduce_ps141 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx141 ^ multm_reduce_mulsc_mulb_pc141;
  assign multm_reduce_ps142 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx142 ^ multm_reduce_mulsc_mulb_pc142;
  assign multm_reduce_ps143 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx143 ^ multm_reduce_mulsc_mulb_pc143;
  assign multm_reduce_ps144 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx144 ^ multm_reduce_mulsc_mulb_pc144;
  assign multm_reduce_ps145 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx145 ^ multm_reduce_mulsc_mulb_pc145;
  assign multm_reduce_ps146 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx146 ^ multm_reduce_mulsc_mulb_pc146;
  assign multm_reduce_ps147 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx147 ^ multm_reduce_mulsc_mulb_pc147;
  assign multm_reduce_ps148 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx148 ^ multm_reduce_mulsc_mulb_pc148;
  assign multm_reduce_ps149 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx149 ^ multm_reduce_mulsc_mulb_pc149;
  assign multm_reduce_ps150 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx150 ^ multm_reduce_mulsc_mulb_pc150;
  assign multm_reduce_ps151 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx151 ^ multm_reduce_mulsc_mulb_pc151;
  assign multm_reduce_ps152 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx152 ^ multm_reduce_mulsc_mulb_pc152;
  assign multm_reduce_ps153 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx153 ^ multm_reduce_mulsc_mulb_pc153;
  assign multm_reduce_ps154 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx154 ^ multm_reduce_mulsc_mulb_pc154;
  assign multm_reduce_ps155 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx155 ^ multm_reduce_mulsc_mulb_pc155;
  assign multm_reduce_ps156 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx156 ^ multm_reduce_mulsc_mulb_pc156;
  assign multm_reduce_ps157 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx157 ^ multm_reduce_mulsc_mulb_pc157;
  assign multm_reduce_ps158 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx158 ^ multm_reduce_mulsc_mulb_pc158;
  assign multm_reduce_ps159 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx159 ^ multm_reduce_mulsc_mulb_pc159;
  assign multm_reduce_ps160 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx160 ^ multm_reduce_mulsc_mulb_pc160;
  assign multm_reduce_ps161 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx161 ^ multm_reduce_mulsc_mulb_pc161;
  assign multm_reduce_ps162 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx162 ^ multm_reduce_mulsc_mulb_pc162;
  assign multm_reduce_ps163 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx163 ^ multm_reduce_mulsc_mulb_pc163;
  assign multm_reduce_ps164 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx164 ^ multm_reduce_mulsc_mulb_pc164;
  assign multm_reduce_ps165 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx165 ^ multm_reduce_mulsc_mulb_pc165;
  assign multm_reduce_ps166 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx166 ^ multm_reduce_mulsc_mulb_pc166;
  assign multm_reduce_ps167 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx167 ^ multm_reduce_mulsc_mulb_pc167;
  assign multm_reduce_ps168 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx168 ^ multm_reduce_mulsc_mulb_pc168;
  assign multm_reduce_ps169 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx169 ^ multm_reduce_mulsc_mulb_pc169;
  assign multm_reduce_ps170 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx170 ^ multm_reduce_mulsc_mulb_pc170;
  assign multm_reduce_ps171 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx171 ^ multm_reduce_mulsc_mulb_pc171;
  assign multm_reduce_ps172 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx172 ^ multm_reduce_mulsc_mulb_pc172;
  assign multm_reduce_ps173 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx173 ^ multm_reduce_mulsc_mulb_pc173;
  assign multm_reduce_ps174 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx174 ^ multm_reduce_mulsc_mulb_pc174;
  assign multm_reduce_ps175 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx175 ^ multm_reduce_mulsc_mulb_pc175;
  assign multm_reduce_ps176 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx176 ^ multm_reduce_mulsc_mulb_pc176;
  assign multm_reduce_ps177 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx177 ^ multm_reduce_mulsc_mulb_pc177;
  assign multm_reduce_ps178 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx178 ^ multm_reduce_mulsc_mulb_pc178;
  assign multm_reduce_ps179 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx179 ^ multm_reduce_mulsc_mulb_pc179;
  assign multm_reduce_ps180 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx180 ^ multm_reduce_mulsc_mulb_pc180;
  assign multm_reduce_ps181 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx181 ^ multm_reduce_mulsc_mulb_pc181;
  assign multm_reduce_ps182 = multm_reduce_mulsc_mulb_add3b1_xor3b_wx182 ^ multm_reduce_mulsc_mulb_pc182;
  assign multm_reduce_ps183 = multm_reduce_mulsc_mulb_add3_xor3_wx ^ multm_reduce_mulsc_mulb_pc183;
  assign multm_reduce_qb = multm_reduce_mulb0_sq0 ^ multm_reduce_sa5;
  assign multm_reduce_qc0 = multm_reduce_mulb0_ps0 & multm_reduce_mulb0_pc0;
  assign multm_reduce_qc1 = multm_reduce_mulb0_ps1 & multm_reduce_mulb0_pc1;
  assign multm_reduce_qc2 = multm_reduce_mulb0_ps2 & multm_reduce_mulb0_pc2;
  assign multm_reduce_qc3 = multm_reduce_mulb0_ps3 & multm_reduce_mulb0_pc3;
  assign multm_reduce_qc4 = multm_reduce_mulb0_ps4 & multm_reduce_mulb0_pc4;
  assign multm_reduce_qc5 = multm_reduce_mulb0_ps5 & multm_reduce_mulb0_pc5;
  assign multm_reduce_qc6 = multm_reduce_mulb0_ps6 & multm_reduce_mulb0_pc6;
  assign multm_reduce_qc7 = multm_reduce_mulb0_ps7 & multm_reduce_mulb0_pc7;
  assign multm_reduce_qc8 = multm_reduce_mulb0_ps8 & multm_reduce_mulb0_pc8;
  assign multm_reduce_qc9 = multm_reduce_mulb0_ps9 & multm_reduce_mulb0_pc9;
  assign multm_reduce_qc10 = multm_reduce_mulb0_ps10 & multm_reduce_mulb0_pc10;
  assign multm_reduce_qc11 = multm_reduce_mulb0_ps11 & multm_reduce_mulb0_pc11;
  assign multm_reduce_qc12 = multm_reduce_mulb0_ps12 & multm_reduce_mulb0_pc12;
  assign multm_reduce_qc13 = multm_reduce_mulb0_ps13 & multm_reduce_mulb0_pc13;
  assign multm_reduce_qc14 = multm_reduce_mulb0_ps14 & multm_reduce_mulb0_pc14;
  assign multm_reduce_qc15 = multm_reduce_mulb0_ps15 & multm_reduce_mulb0_pc15;
  assign multm_reduce_qc16 = multm_reduce_mulb0_ps16 & multm_reduce_mulb0_pc16;
  assign multm_reduce_qc17 = multm_reduce_mulb0_ps17 & multm_reduce_mulb0_pc17;
  assign multm_reduce_qc18 = multm_reduce_mulb0_ps18 & multm_reduce_mulb0_pc18;
  assign multm_reduce_qc19 = multm_reduce_mulb0_ps19 & multm_reduce_mulb0_pc19;
  assign multm_reduce_qc20 = multm_reduce_mulb0_ps20 & multm_reduce_mulb0_pc20;
  assign multm_reduce_qc21 = multm_reduce_mulb0_ps21 & multm_reduce_mulb0_pc21;
  assign multm_reduce_qc22 = multm_reduce_mulb0_ps22 & multm_reduce_mulb0_pc22;
  assign multm_reduce_qc23 = multm_reduce_mulb0_ps23 & multm_reduce_mulb0_pc23;
  assign multm_reduce_qc24 = multm_reduce_mulb0_ps24 & multm_reduce_mulb0_pc24;
  assign multm_reduce_qc25 = multm_reduce_mulb0_ps25 & multm_reduce_mulb0_pc25;
  assign multm_reduce_qc26 = multm_reduce_mulb0_ps26 & multm_reduce_mulb0_pc26;
  assign multm_reduce_qc27 = multm_reduce_mulb0_ps27 & multm_reduce_mulb0_pc27;
  assign multm_reduce_qc28 = multm_reduce_mulb0_ps28 & multm_reduce_mulb0_pc28;
  assign multm_reduce_qc29 = multm_reduce_mulb0_ps29 & multm_reduce_mulb0_pc29;
  assign multm_reduce_qc30 = multm_reduce_mulb0_ps30 & multm_reduce_mulb0_pc30;
  assign multm_reduce_qc31 = multm_reduce_mulb0_ps31 & multm_reduce_mulb0_pc31;
  assign multm_reduce_qc32 = multm_reduce_mulb0_ps32 & multm_reduce_mulb0_pc32;
  assign multm_reduce_qc33 = multm_reduce_mulb0_ps33 & multm_reduce_mulb0_pc33;
  assign multm_reduce_qc34 = multm_reduce_mulb0_ps34 & multm_reduce_mulb0_pc34;
  assign multm_reduce_qc35 = multm_reduce_mulb0_ps35 & multm_reduce_mulb0_pc35;
  assign multm_reduce_qc36 = multm_reduce_mulb0_ps36 & multm_reduce_mulb0_pc36;
  assign multm_reduce_qc37 = multm_reduce_mulb0_ps37 & multm_reduce_mulb0_pc37;
  assign multm_reduce_qc38 = multm_reduce_mulb0_ps38 & multm_reduce_mulb0_pc38;
  assign multm_reduce_qc39 = multm_reduce_mulb0_ps39 & multm_reduce_mulb0_pc39;
  assign multm_reduce_qc40 = multm_reduce_mulb0_ps40 & multm_reduce_mulb0_pc40;
  assign multm_reduce_qc41 = multm_reduce_mulb0_ps41 & multm_reduce_mulb0_pc41;
  assign multm_reduce_qc42 = multm_reduce_mulb0_ps42 & multm_reduce_mulb0_pc42;
  assign multm_reduce_qc43 = multm_reduce_mulb0_ps43 & multm_reduce_mulb0_pc43;
  assign multm_reduce_qc44 = multm_reduce_mulb0_ps44 & multm_reduce_mulb0_pc44;
  assign multm_reduce_qc45 = multm_reduce_mulb0_ps45 & multm_reduce_mulb0_pc45;
  assign multm_reduce_qc46 = multm_reduce_mulb0_ps46 & multm_reduce_mulb0_pc46;
  assign multm_reduce_qc47 = multm_reduce_mulb0_ps47 & multm_reduce_mulb0_pc47;
  assign multm_reduce_qc48 = multm_reduce_mulb0_ps48 & multm_reduce_mulb0_pc48;
  assign multm_reduce_qc49 = multm_reduce_mulb0_ps49 & multm_reduce_mulb0_pc49;
  assign multm_reduce_qc50 = multm_reduce_mulb0_ps50 & multm_reduce_mulb0_pc50;
  assign multm_reduce_qc51 = multm_reduce_mulb0_ps51 & multm_reduce_mulb0_pc51;
  assign multm_reduce_qc52 = multm_reduce_mulb0_ps52 & multm_reduce_mulb0_pc52;
  assign multm_reduce_qc53 = multm_reduce_mulb0_ps53 & multm_reduce_mulb0_pc53;
  assign multm_reduce_qc54 = multm_reduce_mulb0_ps54 & multm_reduce_mulb0_pc54;
  assign multm_reduce_qc55 = multm_reduce_mulb0_ps55 & multm_reduce_mulb0_pc55;
  assign multm_reduce_qc56 = multm_reduce_mulb0_ps56 & multm_reduce_mulb0_pc56;
  assign multm_reduce_qc57 = multm_reduce_mulb0_ps57 & multm_reduce_mulb0_pc57;
  assign multm_reduce_qc58 = multm_reduce_mulb0_ps58 & multm_reduce_mulb0_pc58;
  assign multm_reduce_qc59 = multm_reduce_mulb0_ps59 & multm_reduce_mulb0_pc59;
  assign multm_reduce_qc60 = multm_reduce_mulb0_ps60 & multm_reduce_mulb0_pc60;
  assign multm_reduce_qc61 = multm_reduce_mulb0_ps61 & multm_reduce_mulb0_pc61;
  assign multm_reduce_qc62 = multm_reduce_mulb0_ps62 & multm_reduce_mulb0_pc62;
  assign multm_reduce_qc63 = multm_reduce_mulb0_ps63 & multm_reduce_mulb0_pc63;
  assign multm_reduce_qc64 = multm_reduce_mulb0_ps64 & multm_reduce_mulb0_pc64;
  assign multm_reduce_qc65 = multm_reduce_mulb0_ps65 & multm_reduce_mulb0_pc65;
  assign multm_reduce_qc66 = multm_reduce_mulb0_ps66 & multm_reduce_mulb0_pc66;
  assign multm_reduce_qc67 = multm_reduce_mulb0_ps67 & multm_reduce_mulb0_pc67;
  assign multm_reduce_qc68 = multm_reduce_mulb0_ps68 & multm_reduce_mulb0_pc68;
  assign multm_reduce_qc69 = multm_reduce_mulb0_ps69 & multm_reduce_mulb0_pc69;
  assign multm_reduce_qc70 = multm_reduce_mulb0_ps70 & multm_reduce_mulb0_pc70;
  assign multm_reduce_qc71 = multm_reduce_mulb0_ps71 & multm_reduce_mulb0_pc71;
  assign multm_reduce_qc72 = multm_reduce_mulb0_ps72 & multm_reduce_mulb0_pc72;
  assign multm_reduce_qc73 = multm_reduce_mulb0_ps73 & multm_reduce_mulb0_pc73;
  assign multm_reduce_qc74 = multm_reduce_mulb0_ps74 & multm_reduce_mulb0_pc74;
  assign multm_reduce_qc75 = multm_reduce_mulb0_ps75 & multm_reduce_mulb0_pc75;
  assign multm_reduce_qc76 = multm_reduce_mulb0_ps76 & multm_reduce_mulb0_pc76;
  assign multm_reduce_qc77 = multm_reduce_mulb0_ps77 & multm_reduce_mulb0_pc77;
  assign multm_reduce_qc78 = multm_reduce_mulb0_ps78 & multm_reduce_mulb0_pc78;
  assign multm_reduce_qc79 = multm_reduce_mulb0_ps79 & multm_reduce_mulb0_pc79;
  assign multm_reduce_qc80 = multm_reduce_mulb0_ps80 & multm_reduce_mulb0_pc80;
  assign multm_reduce_qc81 = multm_reduce_mulb0_ps81 & multm_reduce_mulb0_pc81;
  assign multm_reduce_qc82 = multm_reduce_mulb0_ps82 & multm_reduce_mulb0_pc82;
  assign multm_reduce_qc83 = multm_reduce_mulb0_ps83 & multm_reduce_mulb0_pc83;
  assign multm_reduce_qc84 = multm_reduce_mulb0_ps84 & multm_reduce_mulb0_pc84;
  assign multm_reduce_qc85 = multm_reduce_mulb0_ps85 & multm_reduce_mulb0_pc85;
  assign multm_reduce_qc86 = multm_reduce_mulb0_ps86 & multm_reduce_mulb0_pc86;
  assign multm_reduce_qc87 = multm_reduce_mulb0_ps87 & multm_reduce_mulb0_pc87;
  assign multm_reduce_qc88 = multm_reduce_mulb0_ps88 & multm_reduce_mulb0_pc88;
  assign multm_reduce_qc89 = multm_reduce_mulb0_ps89 & multm_reduce_mulb0_pc89;
  assign multm_reduce_qc90 = multm_reduce_mulb0_ps90 & multm_reduce_mulb0_pc90;
  assign multm_reduce_qc91 = multm_reduce_mulb0_ps91 & multm_reduce_mulb0_pc91;
  assign multm_reduce_qc92 = multm_reduce_mulb0_ps92 & multm_reduce_mulb0_pc92;
  assign multm_reduce_qc93 = multm_reduce_mulb0_ps93 & multm_reduce_mulb0_pc93;
  assign multm_reduce_qc94 = multm_reduce_mulb0_ps94 & multm_reduce_mulb0_pc94;
  assign multm_reduce_qc95 = multm_reduce_mulb0_ps95 & multm_reduce_mulb0_pc95;
  assign multm_reduce_qc96 = multm_reduce_mulb0_ps96 & multm_reduce_mulb0_pc96;
  assign multm_reduce_qc97 = multm_reduce_mulb0_ps97 & multm_reduce_mulb0_pc97;
  assign multm_reduce_qc98 = multm_reduce_mulb0_ps98 & multm_reduce_mulb0_pc98;
  assign multm_reduce_qc99 = multm_reduce_mulb0_ps99 & multm_reduce_mulb0_pc99;
  assign multm_reduce_qc100 = multm_reduce_mulb0_ps100 & multm_reduce_mulb0_pc100;
  assign multm_reduce_qc101 = multm_reduce_mulb0_ps101 & multm_reduce_mulb0_pc101;
  assign multm_reduce_qc102 = multm_reduce_mulb0_ps102 & multm_reduce_mulb0_pc102;
  assign multm_reduce_qc103 = multm_reduce_mulb0_ps103 & multm_reduce_mulb0_pc103;
  assign multm_reduce_qc104 = multm_reduce_mulb0_ps104 & multm_reduce_mulb0_pc104;
  assign multm_reduce_qc105 = multm_reduce_mulb0_ps105 & multm_reduce_mulb0_pc105;
  assign multm_reduce_qc106 = multm_reduce_mulb0_ps106 & multm_reduce_mulb0_pc106;
  assign multm_reduce_qc107 = multm_reduce_mulb0_ps107 & multm_reduce_mulb0_pc107;
  assign multm_reduce_qc108 = multm_reduce_mulb0_ps108 & multm_reduce_mulb0_pc108;
  assign multm_reduce_qc109 = multm_reduce_mulb0_ps109 & multm_reduce_mulb0_pc109;
  assign multm_reduce_qc110 = multm_reduce_mulb0_ps110 & multm_reduce_mulb0_pc110;
  assign multm_reduce_qc111 = multm_reduce_mulb0_ps111 & multm_reduce_mulb0_pc111;
  assign multm_reduce_qc112 = multm_reduce_mulb0_ps112 & multm_reduce_mulb0_pc112;
  assign multm_reduce_qc113 = multm_reduce_mulb0_ps113 & multm_reduce_mulb0_pc113;
  assign multm_reduce_qc114 = multm_reduce_mulb0_ps114 & multm_reduce_mulb0_pc114;
  assign multm_reduce_qc115 = multm_reduce_mulb0_ps115 & multm_reduce_mulb0_pc115;
  assign multm_reduce_qc116 = multm_reduce_mulb0_ps116 & multm_reduce_mulb0_pc116;
  assign multm_reduce_qc117 = multm_reduce_mulb0_ps117 & multm_reduce_mulb0_pc117;
  assign multm_reduce_qc118 = multm_reduce_mulb0_ps118 & multm_reduce_mulb0_pc118;
  assign multm_reduce_qc119 = multm_reduce_mulb0_ps119 & multm_reduce_mulb0_pc119;
  assign multm_reduce_qc120 = multm_reduce_mulb0_ps120 & multm_reduce_mulb0_pc120;
  assign multm_reduce_qc121 = multm_reduce_mulb0_ps121 & multm_reduce_mulb0_pc121;
  assign multm_reduce_qc122 = multm_reduce_mulb0_ps122 & multm_reduce_mulb0_pc122;
  assign multm_reduce_qc123 = multm_reduce_mulb0_ps123 & multm_reduce_mulb0_pc123;
  assign multm_reduce_qc124 = multm_reduce_mulb0_ps124 & multm_reduce_mulb0_pc124;
  assign multm_reduce_qc125 = multm_reduce_mulb0_ps125 & multm_reduce_mulb0_pc125;
  assign multm_reduce_qc126 = multm_reduce_mulb0_ps126 & multm_reduce_mulb0_pc126;
  assign multm_reduce_qc127 = multm_reduce_mulb0_ps127 & multm_reduce_mulb0_pc127;
  assign multm_reduce_qc128 = multm_reduce_mulb0_ps128 & multm_reduce_mulb0_pc128;
  assign multm_reduce_qc129 = multm_reduce_mulb0_ps129 & multm_reduce_mulb0_pc129;
  assign multm_reduce_qc130 = multm_reduce_mulb0_ps130 & multm_reduce_mulb0_pc130;
  assign multm_reduce_qc131 = multm_reduce_mulb0_ps131 & multm_reduce_mulb0_pc131;
  assign multm_reduce_qc132 = multm_reduce_mulb0_ps132 & multm_reduce_mulb0_pc132;
  assign multm_reduce_qc133 = multm_reduce_mulb0_ps133 & multm_reduce_mulb0_pc133;
  assign multm_reduce_qc134 = multm_reduce_mulb0_ps134 & multm_reduce_mulb0_pc134;
  assign multm_reduce_qc135 = multm_reduce_mulb0_ps135 & multm_reduce_mulb0_pc135;
  assign multm_reduce_qc136 = multm_reduce_mulb0_ps136 & multm_reduce_mulb0_pc136;
  assign multm_reduce_qc137 = multm_reduce_mulb0_ps137 & multm_reduce_mulb0_pc137;
  assign multm_reduce_qc138 = multm_reduce_mulb0_ps138 & multm_reduce_mulb0_pc138;
  assign multm_reduce_qc139 = multm_reduce_mulb0_ps139 & multm_reduce_mulb0_pc139;
  assign multm_reduce_qc140 = multm_reduce_mulb0_ps140 & multm_reduce_mulb0_pc140;
  assign multm_reduce_qc141 = multm_reduce_mulb0_ps141 & multm_reduce_mulb0_pc141;
  assign multm_reduce_qc142 = multm_reduce_mulb0_ps142 & multm_reduce_mulb0_pc142;
  assign multm_reduce_qc143 = multm_reduce_mulb0_ps143 & multm_reduce_mulb0_pc143;
  assign multm_reduce_qc144 = multm_reduce_mulb0_ps144 & multm_reduce_mulb0_pc144;
  assign multm_reduce_qc145 = multm_reduce_mulb0_ps145 & multm_reduce_mulb0_pc145;
  assign multm_reduce_qc146 = multm_reduce_mulb0_ps146 & multm_reduce_mulb0_pc146;
  assign multm_reduce_qc147 = multm_reduce_mulb0_ps147 & multm_reduce_mulb0_pc147;
  assign multm_reduce_qc148 = multm_reduce_mulb0_ps148 & multm_reduce_mulb0_pc148;
  assign multm_reduce_qc149 = multm_reduce_mulb0_ps149 & multm_reduce_mulb0_pc149;
  assign multm_reduce_qc150 = multm_reduce_mulb0_ps150 & multm_reduce_mulb0_pc150;
  assign multm_reduce_qc151 = multm_reduce_mulb0_ps151 & multm_reduce_mulb0_pc151;
  assign multm_reduce_qc152 = multm_reduce_mulb0_ps152 & multm_reduce_mulb0_pc152;
  assign multm_reduce_qc153 = multm_reduce_mulb0_ps153 & multm_reduce_mulb0_pc153;
  assign multm_reduce_qc154 = multm_reduce_mulb0_ps154 & multm_reduce_mulb0_pc154;
  assign multm_reduce_qc155 = multm_reduce_mulb0_ps155 & multm_reduce_mulb0_pc155;
  assign multm_reduce_qc156 = multm_reduce_mulb0_ps156 & multm_reduce_mulb0_pc156;
  assign multm_reduce_qc157 = multm_reduce_mulb0_ps157 & multm_reduce_mulb0_pc157;
  assign multm_reduce_qc158 = multm_reduce_mulb0_ps158 & multm_reduce_mulb0_pc158;
  assign multm_reduce_qc159 = multm_reduce_mulb0_ps159 & multm_reduce_mulb0_pc159;
  assign multm_reduce_qc160 = multm_reduce_mulb0_ps160 & multm_reduce_mulb0_pc160;
  assign multm_reduce_qc161 = multm_reduce_mulb0_ps161 & multm_reduce_mulb0_pc161;
  assign multm_reduce_qc162 = multm_reduce_mulb0_ps162 & multm_reduce_mulb0_pc162;
  assign multm_reduce_qc163 = multm_reduce_mulb0_ps163 & multm_reduce_mulb0_pc163;
  assign multm_reduce_qc164 = multm_reduce_mulb0_ps164 & multm_reduce_mulb0_pc164;
  assign multm_reduce_qc165 = multm_reduce_mulb0_ps165 & multm_reduce_mulb0_pc165;
  assign multm_reduce_qc166 = multm_reduce_mulb0_ps166 & multm_reduce_mulb0_pc166;
  assign multm_reduce_qc167 = multm_reduce_mulb0_ps167 & multm_reduce_mulb0_pc167;
  assign multm_reduce_qc168 = multm_reduce_mulb0_ps168 & multm_reduce_mulb0_pc168;
  assign multm_reduce_qc169 = multm_reduce_mulb0_ps169 & multm_reduce_mulb0_pc169;
  assign multm_reduce_qc170 = multm_reduce_mulb0_ps170 & multm_reduce_mulb0_pc170;
  assign multm_reduce_qc171 = multm_reduce_mulb0_ps171 & multm_reduce_mulb0_pc171;
  assign multm_reduce_qc172 = multm_reduce_mulb0_ps172 & multm_reduce_mulb0_pc172;
  assign multm_reduce_qc173 = multm_reduce_mulb0_ps173 & multm_reduce_mulb0_pc173;
  assign multm_reduce_qc174 = multm_reduce_mulb0_ps174 & multm_reduce_mulb0_pc174;
  assign multm_reduce_qc175 = multm_reduce_mulb0_ps175 & multm_reduce_mulb0_pc175;
  assign multm_reduce_qc176 = multm_reduce_mulb0_ps176 & multm_reduce_mulb0_pc176;
  assign multm_reduce_qc177 = multm_reduce_mulb0_ps177 & multm_reduce_mulb0_pc177;
  assign multm_reduce_qc178 = multm_reduce_mulb0_ps178 & multm_reduce_mulb0_pc178;
  assign multm_reduce_qc179 = multm_reduce_mulb0_ps179 & multm_reduce_mulb0_pc179;
  assign multm_reduce_qc180 = multm_reduce_mulb0_ps180 & multm_reduce_mulb0_pc180;
  assign multm_reduce_qc181 = multm_reduce_mulb0_ps181 & multm_reduce_mulb0_pc181;
  assign multm_reduce_qc182 = multm_reduce_mulb0_ps182 & multm_reduce_mulb0_pc182;
  assign multm_reduce_qc183 = multm_reduce_mulb0_ps183 & multm_reduce_mulb0_pc183;
  assign multm_reduce_qc184 = multm_reduce_mulb0_add3_maj3_or3_wx | multm_reduce_mulb0_add3_maj3_xy;
  assign multm_reduce_qs0 = multm_reduce_mulb0_ps0 ^ multm_reduce_mulb0_pc0;
  assign multm_reduce_qs1 = multm_reduce_mulb0_ps1 ^ multm_reduce_mulb0_pc1;
  assign multm_reduce_qs2 = multm_reduce_mulb0_ps2 ^ multm_reduce_mulb0_pc2;
  assign multm_reduce_qs3 = multm_reduce_mulb0_ps3 ^ multm_reduce_mulb0_pc3;
  assign multm_reduce_qs4 = multm_reduce_mulb0_ps4 ^ multm_reduce_mulb0_pc4;
  assign multm_reduce_qs5 = multm_reduce_mulb0_ps5 ^ multm_reduce_mulb0_pc5;
  assign multm_reduce_qs6 = multm_reduce_mulb0_ps6 ^ multm_reduce_mulb0_pc6;
  assign multm_reduce_qs7 = multm_reduce_mulb0_ps7 ^ multm_reduce_mulb0_pc7;
  assign multm_reduce_qs8 = multm_reduce_mulb0_ps8 ^ multm_reduce_mulb0_pc8;
  assign multm_reduce_qs9 = multm_reduce_mulb0_ps9 ^ multm_reduce_mulb0_pc9;
  assign multm_reduce_qs10 = multm_reduce_mulb0_ps10 ^ multm_reduce_mulb0_pc10;
  assign multm_reduce_qs11 = multm_reduce_mulb0_ps11 ^ multm_reduce_mulb0_pc11;
  assign multm_reduce_qs12 = multm_reduce_mulb0_ps12 ^ multm_reduce_mulb0_pc12;
  assign multm_reduce_qs13 = multm_reduce_mulb0_ps13 ^ multm_reduce_mulb0_pc13;
  assign multm_reduce_qs14 = multm_reduce_mulb0_ps14 ^ multm_reduce_mulb0_pc14;
  assign multm_reduce_qs15 = multm_reduce_mulb0_ps15 ^ multm_reduce_mulb0_pc15;
  assign multm_reduce_qs16 = multm_reduce_mulb0_ps16 ^ multm_reduce_mulb0_pc16;
  assign multm_reduce_qs17 = multm_reduce_mulb0_ps17 ^ multm_reduce_mulb0_pc17;
  assign multm_reduce_qs18 = multm_reduce_mulb0_ps18 ^ multm_reduce_mulb0_pc18;
  assign multm_reduce_qs19 = multm_reduce_mulb0_ps19 ^ multm_reduce_mulb0_pc19;
  assign multm_reduce_qs20 = multm_reduce_mulb0_ps20 ^ multm_reduce_mulb0_pc20;
  assign multm_reduce_qs21 = multm_reduce_mulb0_ps21 ^ multm_reduce_mulb0_pc21;
  assign multm_reduce_qs22 = multm_reduce_mulb0_ps22 ^ multm_reduce_mulb0_pc22;
  assign multm_reduce_qs23 = multm_reduce_mulb0_ps23 ^ multm_reduce_mulb0_pc23;
  assign multm_reduce_qs24 = multm_reduce_mulb0_ps24 ^ multm_reduce_mulb0_pc24;
  assign multm_reduce_qs25 = multm_reduce_mulb0_ps25 ^ multm_reduce_mulb0_pc25;
  assign multm_reduce_qs26 = multm_reduce_mulb0_ps26 ^ multm_reduce_mulb0_pc26;
  assign multm_reduce_qs27 = multm_reduce_mulb0_ps27 ^ multm_reduce_mulb0_pc27;
  assign multm_reduce_qs28 = multm_reduce_mulb0_ps28 ^ multm_reduce_mulb0_pc28;
  assign multm_reduce_qs29 = multm_reduce_mulb0_ps29 ^ multm_reduce_mulb0_pc29;
  assign multm_reduce_qs30 = multm_reduce_mulb0_ps30 ^ multm_reduce_mulb0_pc30;
  assign multm_reduce_qs31 = multm_reduce_mulb0_ps31 ^ multm_reduce_mulb0_pc31;
  assign multm_reduce_qs32 = multm_reduce_mulb0_ps32 ^ multm_reduce_mulb0_pc32;
  assign multm_reduce_qs33 = multm_reduce_mulb0_ps33 ^ multm_reduce_mulb0_pc33;
  assign multm_reduce_qs34 = multm_reduce_mulb0_ps34 ^ multm_reduce_mulb0_pc34;
  assign multm_reduce_qs35 = multm_reduce_mulb0_ps35 ^ multm_reduce_mulb0_pc35;
  assign multm_reduce_qs36 = multm_reduce_mulb0_ps36 ^ multm_reduce_mulb0_pc36;
  assign multm_reduce_qs37 = multm_reduce_mulb0_ps37 ^ multm_reduce_mulb0_pc37;
  assign multm_reduce_qs38 = multm_reduce_mulb0_ps38 ^ multm_reduce_mulb0_pc38;
  assign multm_reduce_qs39 = multm_reduce_mulb0_ps39 ^ multm_reduce_mulb0_pc39;
  assign multm_reduce_qs40 = multm_reduce_mulb0_ps40 ^ multm_reduce_mulb0_pc40;
  assign multm_reduce_qs41 = multm_reduce_mulb0_ps41 ^ multm_reduce_mulb0_pc41;
  assign multm_reduce_qs42 = multm_reduce_mulb0_ps42 ^ multm_reduce_mulb0_pc42;
  assign multm_reduce_qs43 = multm_reduce_mulb0_ps43 ^ multm_reduce_mulb0_pc43;
  assign multm_reduce_qs44 = multm_reduce_mulb0_ps44 ^ multm_reduce_mulb0_pc44;
  assign multm_reduce_qs45 = multm_reduce_mulb0_ps45 ^ multm_reduce_mulb0_pc45;
  assign multm_reduce_qs46 = multm_reduce_mulb0_ps46 ^ multm_reduce_mulb0_pc46;
  assign multm_reduce_qs47 = multm_reduce_mulb0_ps47 ^ multm_reduce_mulb0_pc47;
  assign multm_reduce_qs48 = multm_reduce_mulb0_ps48 ^ multm_reduce_mulb0_pc48;
  assign multm_reduce_qs49 = multm_reduce_mulb0_ps49 ^ multm_reduce_mulb0_pc49;
  assign multm_reduce_qs50 = multm_reduce_mulb0_ps50 ^ multm_reduce_mulb0_pc50;
  assign multm_reduce_qs51 = multm_reduce_mulb0_ps51 ^ multm_reduce_mulb0_pc51;
  assign multm_reduce_qs52 = multm_reduce_mulb0_ps52 ^ multm_reduce_mulb0_pc52;
  assign multm_reduce_qs53 = multm_reduce_mulb0_ps53 ^ multm_reduce_mulb0_pc53;
  assign multm_reduce_qs54 = multm_reduce_mulb0_ps54 ^ multm_reduce_mulb0_pc54;
  assign multm_reduce_qs55 = multm_reduce_mulb0_ps55 ^ multm_reduce_mulb0_pc55;
  assign multm_reduce_qs56 = multm_reduce_mulb0_ps56 ^ multm_reduce_mulb0_pc56;
  assign multm_reduce_qs57 = multm_reduce_mulb0_ps57 ^ multm_reduce_mulb0_pc57;
  assign multm_reduce_qs58 = multm_reduce_mulb0_ps58 ^ multm_reduce_mulb0_pc58;
  assign multm_reduce_qs59 = multm_reduce_mulb0_ps59 ^ multm_reduce_mulb0_pc59;
  assign multm_reduce_qs60 = multm_reduce_mulb0_ps60 ^ multm_reduce_mulb0_pc60;
  assign multm_reduce_qs61 = multm_reduce_mulb0_ps61 ^ multm_reduce_mulb0_pc61;
  assign multm_reduce_qs62 = multm_reduce_mulb0_ps62 ^ multm_reduce_mulb0_pc62;
  assign multm_reduce_qs63 = multm_reduce_mulb0_ps63 ^ multm_reduce_mulb0_pc63;
  assign multm_reduce_qs64 = multm_reduce_mulb0_ps64 ^ multm_reduce_mulb0_pc64;
  assign multm_reduce_qs65 = multm_reduce_mulb0_ps65 ^ multm_reduce_mulb0_pc65;
  assign multm_reduce_qs66 = multm_reduce_mulb0_ps66 ^ multm_reduce_mulb0_pc66;
  assign multm_reduce_qs67 = multm_reduce_mulb0_ps67 ^ multm_reduce_mulb0_pc67;
  assign multm_reduce_qs68 = multm_reduce_mulb0_ps68 ^ multm_reduce_mulb0_pc68;
  assign multm_reduce_qs69 = multm_reduce_mulb0_ps69 ^ multm_reduce_mulb0_pc69;
  assign multm_reduce_qs70 = multm_reduce_mulb0_ps70 ^ multm_reduce_mulb0_pc70;
  assign multm_reduce_qs71 = multm_reduce_mulb0_ps71 ^ multm_reduce_mulb0_pc71;
  assign multm_reduce_qs72 = multm_reduce_mulb0_ps72 ^ multm_reduce_mulb0_pc72;
  assign multm_reduce_qs73 = multm_reduce_mulb0_ps73 ^ multm_reduce_mulb0_pc73;
  assign multm_reduce_qs74 = multm_reduce_mulb0_ps74 ^ multm_reduce_mulb0_pc74;
  assign multm_reduce_qs75 = multm_reduce_mulb0_ps75 ^ multm_reduce_mulb0_pc75;
  assign multm_reduce_qs76 = multm_reduce_mulb0_ps76 ^ multm_reduce_mulb0_pc76;
  assign multm_reduce_qs77 = multm_reduce_mulb0_ps77 ^ multm_reduce_mulb0_pc77;
  assign multm_reduce_qs78 = multm_reduce_mulb0_ps78 ^ multm_reduce_mulb0_pc78;
  assign multm_reduce_qs79 = multm_reduce_mulb0_ps79 ^ multm_reduce_mulb0_pc79;
  assign multm_reduce_qs80 = multm_reduce_mulb0_ps80 ^ multm_reduce_mulb0_pc80;
  assign multm_reduce_qs81 = multm_reduce_mulb0_ps81 ^ multm_reduce_mulb0_pc81;
  assign multm_reduce_qs82 = multm_reduce_mulb0_ps82 ^ multm_reduce_mulb0_pc82;
  assign multm_reduce_qs83 = multm_reduce_mulb0_ps83 ^ multm_reduce_mulb0_pc83;
  assign multm_reduce_qs84 = multm_reduce_mulb0_ps84 ^ multm_reduce_mulb0_pc84;
  assign multm_reduce_qs85 = multm_reduce_mulb0_ps85 ^ multm_reduce_mulb0_pc85;
  assign multm_reduce_qs86 = multm_reduce_mulb0_ps86 ^ multm_reduce_mulb0_pc86;
  assign multm_reduce_qs87 = multm_reduce_mulb0_ps87 ^ multm_reduce_mulb0_pc87;
  assign multm_reduce_qs88 = multm_reduce_mulb0_ps88 ^ multm_reduce_mulb0_pc88;
  assign multm_reduce_qs89 = multm_reduce_mulb0_ps89 ^ multm_reduce_mulb0_pc89;
  assign multm_reduce_qs90 = multm_reduce_mulb0_ps90 ^ multm_reduce_mulb0_pc90;
  assign multm_reduce_qs91 = multm_reduce_mulb0_ps91 ^ multm_reduce_mulb0_pc91;
  assign multm_reduce_qs92 = multm_reduce_mulb0_ps92 ^ multm_reduce_mulb0_pc92;
  assign multm_reduce_qs93 = multm_reduce_mulb0_ps93 ^ multm_reduce_mulb0_pc93;
  assign multm_reduce_qs94 = multm_reduce_mulb0_ps94 ^ multm_reduce_mulb0_pc94;
  assign multm_reduce_qs95 = multm_reduce_mulb0_ps95 ^ multm_reduce_mulb0_pc95;
  assign multm_reduce_qs96 = multm_reduce_mulb0_ps96 ^ multm_reduce_mulb0_pc96;
  assign multm_reduce_qs97 = multm_reduce_mulb0_ps97 ^ multm_reduce_mulb0_pc97;
  assign multm_reduce_qs98 = multm_reduce_mulb0_ps98 ^ multm_reduce_mulb0_pc98;
  assign multm_reduce_qs99 = multm_reduce_mulb0_ps99 ^ multm_reduce_mulb0_pc99;
  assign multm_reduce_qs100 = multm_reduce_mulb0_ps100 ^ multm_reduce_mulb0_pc100;
  assign multm_reduce_qs101 = multm_reduce_mulb0_ps101 ^ multm_reduce_mulb0_pc101;
  assign multm_reduce_qs102 = multm_reduce_mulb0_ps102 ^ multm_reduce_mulb0_pc102;
  assign multm_reduce_qs103 = multm_reduce_mulb0_ps103 ^ multm_reduce_mulb0_pc103;
  assign multm_reduce_qs104 = multm_reduce_mulb0_ps104 ^ multm_reduce_mulb0_pc104;
  assign multm_reduce_qs105 = multm_reduce_mulb0_ps105 ^ multm_reduce_mulb0_pc105;
  assign multm_reduce_qs106 = multm_reduce_mulb0_ps106 ^ multm_reduce_mulb0_pc106;
  assign multm_reduce_qs107 = multm_reduce_mulb0_ps107 ^ multm_reduce_mulb0_pc107;
  assign multm_reduce_qs108 = multm_reduce_mulb0_ps108 ^ multm_reduce_mulb0_pc108;
  assign multm_reduce_qs109 = multm_reduce_mulb0_ps109 ^ multm_reduce_mulb0_pc109;
  assign multm_reduce_qs110 = multm_reduce_mulb0_ps110 ^ multm_reduce_mulb0_pc110;
  assign multm_reduce_qs111 = multm_reduce_mulb0_ps111 ^ multm_reduce_mulb0_pc111;
  assign multm_reduce_qs112 = multm_reduce_mulb0_ps112 ^ multm_reduce_mulb0_pc112;
  assign multm_reduce_qs113 = multm_reduce_mulb0_ps113 ^ multm_reduce_mulb0_pc113;
  assign multm_reduce_qs114 = multm_reduce_mulb0_ps114 ^ multm_reduce_mulb0_pc114;
  assign multm_reduce_qs115 = multm_reduce_mulb0_ps115 ^ multm_reduce_mulb0_pc115;
  assign multm_reduce_qs116 = multm_reduce_mulb0_ps116 ^ multm_reduce_mulb0_pc116;
  assign multm_reduce_qs117 = multm_reduce_mulb0_ps117 ^ multm_reduce_mulb0_pc117;
  assign multm_reduce_qs118 = multm_reduce_mulb0_ps118 ^ multm_reduce_mulb0_pc118;
  assign multm_reduce_qs119 = multm_reduce_mulb0_ps119 ^ multm_reduce_mulb0_pc119;
  assign multm_reduce_qs120 = multm_reduce_mulb0_ps120 ^ multm_reduce_mulb0_pc120;
  assign multm_reduce_qs121 = multm_reduce_mulb0_ps121 ^ multm_reduce_mulb0_pc121;
  assign multm_reduce_qs122 = multm_reduce_mulb0_ps122 ^ multm_reduce_mulb0_pc122;
  assign multm_reduce_qs123 = multm_reduce_mulb0_ps123 ^ multm_reduce_mulb0_pc123;
  assign multm_reduce_qs124 = multm_reduce_mulb0_ps124 ^ multm_reduce_mulb0_pc124;
  assign multm_reduce_qs125 = multm_reduce_mulb0_ps125 ^ multm_reduce_mulb0_pc125;
  assign multm_reduce_qs126 = multm_reduce_mulb0_ps126 ^ multm_reduce_mulb0_pc126;
  assign multm_reduce_qs127 = multm_reduce_mulb0_ps127 ^ multm_reduce_mulb0_pc127;
  assign multm_reduce_qs128 = multm_reduce_mulb0_ps128 ^ multm_reduce_mulb0_pc128;
  assign multm_reduce_qs129 = multm_reduce_mulb0_ps129 ^ multm_reduce_mulb0_pc129;
  assign multm_reduce_qs130 = multm_reduce_mulb0_ps130 ^ multm_reduce_mulb0_pc130;
  assign multm_reduce_qs131 = multm_reduce_mulb0_ps131 ^ multm_reduce_mulb0_pc131;
  assign multm_reduce_qs132 = multm_reduce_mulb0_ps132 ^ multm_reduce_mulb0_pc132;
  assign multm_reduce_qs133 = multm_reduce_mulb0_ps133 ^ multm_reduce_mulb0_pc133;
  assign multm_reduce_qs134 = multm_reduce_mulb0_ps134 ^ multm_reduce_mulb0_pc134;
  assign multm_reduce_qs135 = multm_reduce_mulb0_ps135 ^ multm_reduce_mulb0_pc135;
  assign multm_reduce_qs136 = multm_reduce_mulb0_ps136 ^ multm_reduce_mulb0_pc136;
  assign multm_reduce_qs137 = multm_reduce_mulb0_ps137 ^ multm_reduce_mulb0_pc137;
  assign multm_reduce_qs138 = multm_reduce_mulb0_ps138 ^ multm_reduce_mulb0_pc138;
  assign multm_reduce_qs139 = multm_reduce_mulb0_ps139 ^ multm_reduce_mulb0_pc139;
  assign multm_reduce_qs140 = multm_reduce_mulb0_ps140 ^ multm_reduce_mulb0_pc140;
  assign multm_reduce_qs141 = multm_reduce_mulb0_ps141 ^ multm_reduce_mulb0_pc141;
  assign multm_reduce_qs142 = multm_reduce_mulb0_ps142 ^ multm_reduce_mulb0_pc142;
  assign multm_reduce_qs143 = multm_reduce_mulb0_ps143 ^ multm_reduce_mulb0_pc143;
  assign multm_reduce_qs144 = multm_reduce_mulb0_ps144 ^ multm_reduce_mulb0_pc144;
  assign multm_reduce_qs145 = multm_reduce_mulb0_ps145 ^ multm_reduce_mulb0_pc145;
  assign multm_reduce_qs146 = multm_reduce_mulb0_ps146 ^ multm_reduce_mulb0_pc146;
  assign multm_reduce_qs147 = multm_reduce_mulb0_ps147 ^ multm_reduce_mulb0_pc147;
  assign multm_reduce_qs148 = multm_reduce_mulb0_ps148 ^ multm_reduce_mulb0_pc148;
  assign multm_reduce_qs149 = multm_reduce_mulb0_ps149 ^ multm_reduce_mulb0_pc149;
  assign multm_reduce_qs150 = multm_reduce_mulb0_ps150 ^ multm_reduce_mulb0_pc150;
  assign multm_reduce_qs151 = multm_reduce_mulb0_ps151 ^ multm_reduce_mulb0_pc151;
  assign multm_reduce_qs152 = multm_reduce_mulb0_ps152 ^ multm_reduce_mulb0_pc152;
  assign multm_reduce_qs153 = multm_reduce_mulb0_ps153 ^ multm_reduce_mulb0_pc153;
  assign multm_reduce_qs154 = multm_reduce_mulb0_ps154 ^ multm_reduce_mulb0_pc154;
  assign multm_reduce_qs155 = multm_reduce_mulb0_ps155 ^ multm_reduce_mulb0_pc155;
  assign multm_reduce_qs156 = multm_reduce_mulb0_ps156 ^ multm_reduce_mulb0_pc156;
  assign multm_reduce_qs157 = multm_reduce_mulb0_ps157 ^ multm_reduce_mulb0_pc157;
  assign multm_reduce_qs158 = multm_reduce_mulb0_ps158 ^ multm_reduce_mulb0_pc158;
  assign multm_reduce_qs159 = multm_reduce_mulb0_ps159 ^ multm_reduce_mulb0_pc159;
  assign multm_reduce_qs160 = multm_reduce_mulb0_ps160 ^ multm_reduce_mulb0_pc160;
  assign multm_reduce_qs161 = multm_reduce_mulb0_ps161 ^ multm_reduce_mulb0_pc161;
  assign multm_reduce_qs162 = multm_reduce_mulb0_ps162 ^ multm_reduce_mulb0_pc162;
  assign multm_reduce_qs163 = multm_reduce_mulb0_ps163 ^ multm_reduce_mulb0_pc163;
  assign multm_reduce_qs164 = multm_reduce_mulb0_ps164 ^ multm_reduce_mulb0_pc164;
  assign multm_reduce_qs165 = multm_reduce_mulb0_ps165 ^ multm_reduce_mulb0_pc165;
  assign multm_reduce_qs166 = multm_reduce_mulb0_ps166 ^ multm_reduce_mulb0_pc166;
  assign multm_reduce_qs167 = multm_reduce_mulb0_ps167 ^ multm_reduce_mulb0_pc167;
  assign multm_reduce_qs168 = multm_reduce_mulb0_ps168 ^ multm_reduce_mulb0_pc168;
  assign multm_reduce_qs169 = multm_reduce_mulb0_ps169 ^ multm_reduce_mulb0_pc169;
  assign multm_reduce_qs170 = multm_reduce_mulb0_ps170 ^ multm_reduce_mulb0_pc170;
  assign multm_reduce_qs171 = multm_reduce_mulb0_ps171 ^ multm_reduce_mulb0_pc171;
  assign multm_reduce_qs172 = multm_reduce_mulb0_ps172 ^ multm_reduce_mulb0_pc172;
  assign multm_reduce_qs173 = multm_reduce_mulb0_ps173 ^ multm_reduce_mulb0_pc173;
  assign multm_reduce_qs174 = multm_reduce_mulb0_ps174 ^ multm_reduce_mulb0_pc174;
  assign multm_reduce_qs175 = multm_reduce_mulb0_ps175 ^ multm_reduce_mulb0_pc175;
  assign multm_reduce_qs176 = multm_reduce_mulb0_ps176 ^ multm_reduce_mulb0_pc176;
  assign multm_reduce_qs177 = multm_reduce_mulb0_ps177 ^ multm_reduce_mulb0_pc177;
  assign multm_reduce_qs178 = multm_reduce_mulb0_ps178 ^ multm_reduce_mulb0_pc178;
  assign multm_reduce_qs179 = multm_reduce_mulb0_ps179 ^ multm_reduce_mulb0_pc179;
  assign multm_reduce_qs180 = multm_reduce_mulb0_ps180 ^ multm_reduce_mulb0_pc180;
  assign multm_reduce_qs181 = multm_reduce_mulb0_ps181 ^ multm_reduce_mulb0_pc181;
  assign multm_reduce_qs182 = multm_reduce_mulb0_ps182 ^ multm_reduce_mulb0_pc182;
  assign multm_reduce_qs183 = multm_reduce_mulb0_ps183 ^ multm_reduce_mulb0_pc183;
  assign multm_reduce_qs184 = multm_reduce_mulb0_add3_xor3_wx ^ multm_reduce_mulb0_pc184;
  assign multm_reduce_sticky_q = xn2 & multm_reduce_sd0;
  assign multm_reduce_vb = multm_reduce_mulb1_sq0 ^ multm_reduce_qb2;
  assign multm_reduce_vc0 = multm_reduce_mulb1_ps0 & multm_reduce_mulb1_pc0;
  assign multm_reduce_vc1 = multm_reduce_mulb1_ps1 & multm_reduce_mulb1_pc1;
  assign multm_reduce_vc2 = multm_reduce_mulb1_ps2 & multm_reduce_mulb1_pc2;
  assign multm_reduce_vc3 = multm_reduce_mulb1_ps3 & multm_reduce_mulb1_pc3;
  assign multm_reduce_vc4 = multm_reduce_mulb1_ps4 & multm_reduce_mulb1_pc4;
  assign multm_reduce_vc5 = multm_reduce_mulb1_ps5 & multm_reduce_mulb1_pc5;
  assign multm_reduce_vc6 = multm_reduce_mulb1_ps6 & multm_reduce_mulb1_pc6;
  assign multm_reduce_vc7 = multm_reduce_mulb1_ps7 & multm_reduce_mulb1_pc7;
  assign multm_reduce_vc8 = multm_reduce_mulb1_ps8 & multm_reduce_mulb1_pc8;
  assign multm_reduce_vc9 = multm_reduce_mulb1_ps9 & multm_reduce_mulb1_pc9;
  assign multm_reduce_vc10 = multm_reduce_mulb1_ps10 & multm_reduce_mulb1_pc10;
  assign multm_reduce_vc11 = multm_reduce_mulb1_ps11 & multm_reduce_mulb1_pc11;
  assign multm_reduce_vc12 = multm_reduce_mulb1_ps12 & multm_reduce_mulb1_pc12;
  assign multm_reduce_vc13 = multm_reduce_mulb1_ps13 & multm_reduce_mulb1_pc13;
  assign multm_reduce_vc14 = multm_reduce_mulb1_ps14 & multm_reduce_mulb1_pc14;
  assign multm_reduce_vc15 = multm_reduce_mulb1_ps15 & multm_reduce_mulb1_pc15;
  assign multm_reduce_vc16 = multm_reduce_mulb1_ps16 & multm_reduce_mulb1_pc16;
  assign multm_reduce_vc17 = multm_reduce_mulb1_ps17 & multm_reduce_mulb1_pc17;
  assign multm_reduce_vc18 = multm_reduce_mulb1_ps18 & multm_reduce_mulb1_pc18;
  assign multm_reduce_vc19 = multm_reduce_mulb1_ps19 & multm_reduce_mulb1_pc19;
  assign multm_reduce_vc20 = multm_reduce_mulb1_ps20 & multm_reduce_mulb1_pc20;
  assign multm_reduce_vc21 = multm_reduce_mulb1_ps21 & multm_reduce_mulb1_pc21;
  assign multm_reduce_vc22 = multm_reduce_mulb1_ps22 & multm_reduce_mulb1_pc22;
  assign multm_reduce_vc23 = multm_reduce_mulb1_ps23 & multm_reduce_mulb1_pc23;
  assign multm_reduce_vc24 = multm_reduce_mulb1_ps24 & multm_reduce_mulb1_pc24;
  assign multm_reduce_vc25 = multm_reduce_mulb1_ps25 & multm_reduce_mulb1_pc25;
  assign multm_reduce_vc26 = multm_reduce_mulb1_ps26 & multm_reduce_mulb1_pc26;
  assign multm_reduce_vc27 = multm_reduce_mulb1_ps27 & multm_reduce_mulb1_pc27;
  assign multm_reduce_vc28 = multm_reduce_mulb1_ps28 & multm_reduce_mulb1_pc28;
  assign multm_reduce_vc29 = multm_reduce_mulb1_ps29 & multm_reduce_mulb1_pc29;
  assign multm_reduce_vc30 = multm_reduce_mulb1_ps30 & multm_reduce_mulb1_pc30;
  assign multm_reduce_vc31 = multm_reduce_mulb1_ps31 & multm_reduce_mulb1_pc31;
  assign multm_reduce_vc32 = multm_reduce_mulb1_ps32 & multm_reduce_mulb1_pc32;
  assign multm_reduce_vc33 = multm_reduce_mulb1_ps33 & multm_reduce_mulb1_pc33;
  assign multm_reduce_vc34 = multm_reduce_mulb1_ps34 & multm_reduce_mulb1_pc34;
  assign multm_reduce_vc35 = multm_reduce_mulb1_ps35 & multm_reduce_mulb1_pc35;
  assign multm_reduce_vc36 = multm_reduce_mulb1_ps36 & multm_reduce_mulb1_pc36;
  assign multm_reduce_vc37 = multm_reduce_mulb1_ps37 & multm_reduce_mulb1_pc37;
  assign multm_reduce_vc38 = multm_reduce_mulb1_ps38 & multm_reduce_mulb1_pc38;
  assign multm_reduce_vc39 = multm_reduce_mulb1_ps39 & multm_reduce_mulb1_pc39;
  assign multm_reduce_vc40 = multm_reduce_mulb1_ps40 & multm_reduce_mulb1_pc40;
  assign multm_reduce_vc41 = multm_reduce_mulb1_ps41 & multm_reduce_mulb1_pc41;
  assign multm_reduce_vc42 = multm_reduce_mulb1_ps42 & multm_reduce_mulb1_pc42;
  assign multm_reduce_vc43 = multm_reduce_mulb1_ps43 & multm_reduce_mulb1_pc43;
  assign multm_reduce_vc44 = multm_reduce_mulb1_ps44 & multm_reduce_mulb1_pc44;
  assign multm_reduce_vc45 = multm_reduce_mulb1_ps45 & multm_reduce_mulb1_pc45;
  assign multm_reduce_vc46 = multm_reduce_mulb1_ps46 & multm_reduce_mulb1_pc46;
  assign multm_reduce_vc47 = multm_reduce_mulb1_ps47 & multm_reduce_mulb1_pc47;
  assign multm_reduce_vc48 = multm_reduce_mulb1_ps48 & multm_reduce_mulb1_pc48;
  assign multm_reduce_vc49 = multm_reduce_mulb1_ps49 & multm_reduce_mulb1_pc49;
  assign multm_reduce_vc50 = multm_reduce_mulb1_ps50 & multm_reduce_mulb1_pc50;
  assign multm_reduce_vc51 = multm_reduce_mulb1_ps51 & multm_reduce_mulb1_pc51;
  assign multm_reduce_vc52 = multm_reduce_mulb1_ps52 & multm_reduce_mulb1_pc52;
  assign multm_reduce_vc53 = multm_reduce_mulb1_ps53 & multm_reduce_mulb1_pc53;
  assign multm_reduce_vc54 = multm_reduce_mulb1_ps54 & multm_reduce_mulb1_pc54;
  assign multm_reduce_vc55 = multm_reduce_mulb1_ps55 & multm_reduce_mulb1_pc55;
  assign multm_reduce_vc56 = multm_reduce_mulb1_ps56 & multm_reduce_mulb1_pc56;
  assign multm_reduce_vc57 = multm_reduce_mulb1_ps57 & multm_reduce_mulb1_pc57;
  assign multm_reduce_vc58 = multm_reduce_mulb1_ps58 & multm_reduce_mulb1_pc58;
  assign multm_reduce_vc59 = multm_reduce_mulb1_ps59 & multm_reduce_mulb1_pc59;
  assign multm_reduce_vc60 = multm_reduce_mulb1_ps60 & multm_reduce_mulb1_pc60;
  assign multm_reduce_vc61 = multm_reduce_mulb1_ps61 & multm_reduce_mulb1_pc61;
  assign multm_reduce_vc62 = multm_reduce_mulb1_ps62 & multm_reduce_mulb1_pc62;
  assign multm_reduce_vc63 = multm_reduce_mulb1_ps63 & multm_reduce_mulb1_pc63;
  assign multm_reduce_vc64 = multm_reduce_mulb1_ps64 & multm_reduce_mulb1_pc64;
  assign multm_reduce_vc65 = multm_reduce_mulb1_ps65 & multm_reduce_mulb1_pc65;
  assign multm_reduce_vc66 = multm_reduce_mulb1_ps66 & multm_reduce_mulb1_pc66;
  assign multm_reduce_vc67 = multm_reduce_mulb1_ps67 & multm_reduce_mulb1_pc67;
  assign multm_reduce_vc68 = multm_reduce_mulb1_ps68 & multm_reduce_mulb1_pc68;
  assign multm_reduce_vc69 = multm_reduce_mulb1_ps69 & multm_reduce_mulb1_pc69;
  assign multm_reduce_vc70 = multm_reduce_mulb1_ps70 & multm_reduce_mulb1_pc70;
  assign multm_reduce_vc71 = multm_reduce_mulb1_ps71 & multm_reduce_mulb1_pc71;
  assign multm_reduce_vc72 = multm_reduce_mulb1_ps72 & multm_reduce_mulb1_pc72;
  assign multm_reduce_vc73 = multm_reduce_mulb1_ps73 & multm_reduce_mulb1_pc73;
  assign multm_reduce_vc74 = multm_reduce_mulb1_ps74 & multm_reduce_mulb1_pc74;
  assign multm_reduce_vc75 = multm_reduce_mulb1_ps75 & multm_reduce_mulb1_pc75;
  assign multm_reduce_vc76 = multm_reduce_mulb1_ps76 & multm_reduce_mulb1_pc76;
  assign multm_reduce_vc77 = multm_reduce_mulb1_ps77 & multm_reduce_mulb1_pc77;
  assign multm_reduce_vc78 = multm_reduce_mulb1_ps78 & multm_reduce_mulb1_pc78;
  assign multm_reduce_vc79 = multm_reduce_mulb1_ps79 & multm_reduce_mulb1_pc79;
  assign multm_reduce_vc80 = multm_reduce_mulb1_ps80 & multm_reduce_mulb1_pc80;
  assign multm_reduce_vc81 = multm_reduce_mulb1_ps81 & multm_reduce_mulb1_pc81;
  assign multm_reduce_vc82 = multm_reduce_mulb1_ps82 & multm_reduce_mulb1_pc82;
  assign multm_reduce_vc83 = multm_reduce_mulb1_ps83 & multm_reduce_mulb1_pc83;
  assign multm_reduce_vc84 = multm_reduce_mulb1_ps84 & multm_reduce_mulb1_pc84;
  assign multm_reduce_vc85 = multm_reduce_mulb1_ps85 & multm_reduce_mulb1_pc85;
  assign multm_reduce_vc86 = multm_reduce_mulb1_ps86 & multm_reduce_mulb1_pc86;
  assign multm_reduce_vc87 = multm_reduce_mulb1_ps87 & multm_reduce_mulb1_pc87;
  assign multm_reduce_vc88 = multm_reduce_mulb1_ps88 & multm_reduce_mulb1_pc88;
  assign multm_reduce_vc89 = multm_reduce_mulb1_ps89 & multm_reduce_mulb1_pc89;
  assign multm_reduce_vc90 = multm_reduce_mulb1_ps90 & multm_reduce_mulb1_pc90;
  assign multm_reduce_vc91 = multm_reduce_mulb1_ps91 & multm_reduce_mulb1_pc91;
  assign multm_reduce_vc92 = multm_reduce_mulb1_ps92 & multm_reduce_mulb1_pc92;
  assign multm_reduce_vc93 = multm_reduce_mulb1_ps93 & multm_reduce_mulb1_pc93;
  assign multm_reduce_vc94 = multm_reduce_mulb1_ps94 & multm_reduce_mulb1_pc94;
  assign multm_reduce_vc95 = multm_reduce_mulb1_ps95 & multm_reduce_mulb1_pc95;
  assign multm_reduce_vc96 = multm_reduce_mulb1_ps96 & multm_reduce_mulb1_pc96;
  assign multm_reduce_vc97 = multm_reduce_mulb1_ps97 & multm_reduce_mulb1_pc97;
  assign multm_reduce_vc98 = multm_reduce_mulb1_ps98 & multm_reduce_mulb1_pc98;
  assign multm_reduce_vc99 = multm_reduce_mulb1_ps99 & multm_reduce_mulb1_pc99;
  assign multm_reduce_vc100 = multm_reduce_mulb1_ps100 & multm_reduce_mulb1_pc100;
  assign multm_reduce_vc101 = multm_reduce_mulb1_ps101 & multm_reduce_mulb1_pc101;
  assign multm_reduce_vc102 = multm_reduce_mulb1_ps102 & multm_reduce_mulb1_pc102;
  assign multm_reduce_vc103 = multm_reduce_mulb1_ps103 & multm_reduce_mulb1_pc103;
  assign multm_reduce_vc104 = multm_reduce_mulb1_ps104 & multm_reduce_mulb1_pc104;
  assign multm_reduce_vc105 = multm_reduce_mulb1_ps105 & multm_reduce_mulb1_pc105;
  assign multm_reduce_vc106 = multm_reduce_mulb1_ps106 & multm_reduce_mulb1_pc106;
  assign multm_reduce_vc107 = multm_reduce_mulb1_ps107 & multm_reduce_mulb1_pc107;
  assign multm_reduce_vc108 = multm_reduce_mulb1_ps108 & multm_reduce_mulb1_pc108;
  assign multm_reduce_vc109 = multm_reduce_mulb1_ps109 & multm_reduce_mulb1_pc109;
  assign multm_reduce_vc110 = multm_reduce_mulb1_ps110 & multm_reduce_mulb1_pc110;
  assign multm_reduce_vc111 = multm_reduce_mulb1_ps111 & multm_reduce_mulb1_pc111;
  assign multm_reduce_vc112 = multm_reduce_mulb1_ps112 & multm_reduce_mulb1_pc112;
  assign multm_reduce_vc113 = multm_reduce_mulb1_ps113 & multm_reduce_mulb1_pc113;
  assign multm_reduce_vc114 = multm_reduce_mulb1_ps114 & multm_reduce_mulb1_pc114;
  assign multm_reduce_vc115 = multm_reduce_mulb1_ps115 & multm_reduce_mulb1_pc115;
  assign multm_reduce_vc116 = multm_reduce_mulb1_ps116 & multm_reduce_mulb1_pc116;
  assign multm_reduce_vc117 = multm_reduce_mulb1_ps117 & multm_reduce_mulb1_pc117;
  assign multm_reduce_vc118 = multm_reduce_mulb1_ps118 & multm_reduce_mulb1_pc118;
  assign multm_reduce_vc119 = multm_reduce_mulb1_ps119 & multm_reduce_mulb1_pc119;
  assign multm_reduce_vc120 = multm_reduce_mulb1_ps120 & multm_reduce_mulb1_pc120;
  assign multm_reduce_vc121 = multm_reduce_mulb1_ps121 & multm_reduce_mulb1_pc121;
  assign multm_reduce_vc122 = multm_reduce_mulb1_ps122 & multm_reduce_mulb1_pc122;
  assign multm_reduce_vc123 = multm_reduce_mulb1_ps123 & multm_reduce_mulb1_pc123;
  assign multm_reduce_vc124 = multm_reduce_mulb1_ps124 & multm_reduce_mulb1_pc124;
  assign multm_reduce_vc125 = multm_reduce_mulb1_ps125 & multm_reduce_mulb1_pc125;
  assign multm_reduce_vc126 = multm_reduce_mulb1_ps126 & multm_reduce_mulb1_pc126;
  assign multm_reduce_vc127 = multm_reduce_mulb1_ps127 & multm_reduce_mulb1_pc127;
  assign multm_reduce_vc128 = multm_reduce_mulb1_ps128 & multm_reduce_mulb1_pc128;
  assign multm_reduce_vc129 = multm_reduce_mulb1_ps129 & multm_reduce_mulb1_pc129;
  assign multm_reduce_vc130 = multm_reduce_mulb1_ps130 & multm_reduce_mulb1_pc130;
  assign multm_reduce_vc131 = multm_reduce_mulb1_ps131 & multm_reduce_mulb1_pc131;
  assign multm_reduce_vc132 = multm_reduce_mulb1_ps132 & multm_reduce_mulb1_pc132;
  assign multm_reduce_vc133 = multm_reduce_mulb1_ps133 & multm_reduce_mulb1_pc133;
  assign multm_reduce_vc134 = multm_reduce_mulb1_ps134 & multm_reduce_mulb1_pc134;
  assign multm_reduce_vc135 = multm_reduce_mulb1_ps135 & multm_reduce_mulb1_pc135;
  assign multm_reduce_vc136 = multm_reduce_mulb1_ps136 & multm_reduce_mulb1_pc136;
  assign multm_reduce_vc137 = multm_reduce_mulb1_ps137 & multm_reduce_mulb1_pc137;
  assign multm_reduce_vc138 = multm_reduce_mulb1_ps138 & multm_reduce_mulb1_pc138;
  assign multm_reduce_vc139 = multm_reduce_mulb1_ps139 & multm_reduce_mulb1_pc139;
  assign multm_reduce_vc140 = multm_reduce_mulb1_ps140 & multm_reduce_mulb1_pc140;
  assign multm_reduce_vc141 = multm_reduce_mulb1_ps141 & multm_reduce_mulb1_pc141;
  assign multm_reduce_vc142 = multm_reduce_mulb1_ps142 & multm_reduce_mulb1_pc142;
  assign multm_reduce_vc143 = multm_reduce_mulb1_ps143 & multm_reduce_mulb1_pc143;
  assign multm_reduce_vc144 = multm_reduce_mulb1_ps144 & multm_reduce_mulb1_pc144;
  assign multm_reduce_vc145 = multm_reduce_mulb1_ps145 & multm_reduce_mulb1_pc145;
  assign multm_reduce_vc146 = multm_reduce_mulb1_ps146 & multm_reduce_mulb1_pc146;
  assign multm_reduce_vc147 = multm_reduce_mulb1_ps147 & multm_reduce_mulb1_pc147;
  assign multm_reduce_vc148 = multm_reduce_mulb1_ps148 & multm_reduce_mulb1_pc148;
  assign multm_reduce_vc149 = multm_reduce_mulb1_ps149 & multm_reduce_mulb1_pc149;
  assign multm_reduce_vc150 = multm_reduce_mulb1_ps150 & multm_reduce_mulb1_pc150;
  assign multm_reduce_vc151 = multm_reduce_mulb1_ps151 & multm_reduce_mulb1_pc151;
  assign multm_reduce_vc152 = multm_reduce_mulb1_ps152 & multm_reduce_mulb1_pc152;
  assign multm_reduce_vc153 = multm_reduce_mulb1_ps153 & multm_reduce_mulb1_pc153;
  assign multm_reduce_vc154 = multm_reduce_mulb1_ps154 & multm_reduce_mulb1_pc154;
  assign multm_reduce_vc155 = multm_reduce_mulb1_ps155 & multm_reduce_mulb1_pc155;
  assign multm_reduce_vc156 = multm_reduce_mulb1_ps156 & multm_reduce_mulb1_pc156;
  assign multm_reduce_vc157 = multm_reduce_mulb1_ps157 & multm_reduce_mulb1_pc157;
  assign multm_reduce_vc158 = multm_reduce_mulb1_ps158 & multm_reduce_mulb1_pc158;
  assign multm_reduce_vc159 = multm_reduce_mulb1_ps159 & multm_reduce_mulb1_pc159;
  assign multm_reduce_vc160 = multm_reduce_mulb1_ps160 & multm_reduce_mulb1_pc160;
  assign multm_reduce_vc161 = multm_reduce_mulb1_ps161 & multm_reduce_mulb1_pc161;
  assign multm_reduce_vc162 = multm_reduce_mulb1_ps162 & multm_reduce_mulb1_pc162;
  assign multm_reduce_vc163 = multm_reduce_mulb1_ps163 & multm_reduce_mulb1_pc163;
  assign multm_reduce_vc164 = multm_reduce_mulb1_ps164 & multm_reduce_mulb1_pc164;
  assign multm_reduce_vc165 = multm_reduce_mulb1_ps165 & multm_reduce_mulb1_pc165;
  assign multm_reduce_vc166 = multm_reduce_mulb1_ps166 & multm_reduce_mulb1_pc166;
  assign multm_reduce_vc167 = multm_reduce_mulb1_ps167 & multm_reduce_mulb1_pc167;
  assign multm_reduce_vc168 = multm_reduce_mulb1_ps168 & multm_reduce_mulb1_pc168;
  assign multm_reduce_vc169 = multm_reduce_mulb1_ps169 & multm_reduce_mulb1_pc169;
  assign multm_reduce_vc170 = multm_reduce_mulb1_ps170 & multm_reduce_mulb1_pc170;
  assign multm_reduce_vc171 = multm_reduce_mulb1_ps171 & multm_reduce_mulb1_pc171;
  assign multm_reduce_vc172 = multm_reduce_mulb1_ps172 & multm_reduce_mulb1_pc172;
  assign multm_reduce_vc173 = multm_reduce_mulb1_ps173 & multm_reduce_mulb1_pc173;
  assign multm_reduce_vc174 = multm_reduce_mulb1_ps174 & multm_reduce_mulb1_pc174;
  assign multm_reduce_vc175 = multm_reduce_mulb1_ps175 & multm_reduce_mulb1_pc175;
  assign multm_reduce_vc176 = multm_reduce_mulb1_ps176 & multm_reduce_mulb1_pc176;
  assign multm_reduce_vc177 = multm_reduce_mulb1_ps177 & multm_reduce_mulb1_pc177;
  assign multm_reduce_vc178 = multm_reduce_mulb1_ps178 & multm_reduce_mulb1_pc178;
  assign multm_reduce_vc179 = multm_reduce_mulb1_ps179 & multm_reduce_mulb1_pc179;
  assign multm_reduce_vc180 = multm_reduce_mulb1_ps180 & multm_reduce_mulb1_pc180;
  assign multm_reduce_vc181 = multm_reduce_mulb1_ps181 & multm_reduce_mulb1_pc181;
  assign multm_reduce_vc182 = multm_reduce_mulb1_add3_maj3_or3_wx | multm_reduce_mulb1_add3_maj3_xy;
  assign multm_reduce_vs0 = multm_reduce_mulb1_ps0 ^ multm_reduce_mulb1_pc0;
  assign multm_reduce_vs1 = multm_reduce_mulb1_ps1 ^ multm_reduce_mulb1_pc1;
  assign multm_reduce_vs2 = multm_reduce_mulb1_ps2 ^ multm_reduce_mulb1_pc2;
  assign multm_reduce_vs3 = multm_reduce_mulb1_ps3 ^ multm_reduce_mulb1_pc3;
  assign multm_reduce_vs4 = multm_reduce_mulb1_ps4 ^ multm_reduce_mulb1_pc4;
  assign multm_reduce_vs5 = multm_reduce_mulb1_ps5 ^ multm_reduce_mulb1_pc5;
  assign multm_reduce_vs6 = multm_reduce_mulb1_ps6 ^ multm_reduce_mulb1_pc6;
  assign multm_reduce_vs7 = multm_reduce_mulb1_ps7 ^ multm_reduce_mulb1_pc7;
  assign multm_reduce_vs8 = multm_reduce_mulb1_ps8 ^ multm_reduce_mulb1_pc8;
  assign multm_reduce_vs9 = multm_reduce_mulb1_ps9 ^ multm_reduce_mulb1_pc9;
  assign multm_reduce_vs10 = multm_reduce_mulb1_ps10 ^ multm_reduce_mulb1_pc10;
  assign multm_reduce_vs11 = multm_reduce_mulb1_ps11 ^ multm_reduce_mulb1_pc11;
  assign multm_reduce_vs12 = multm_reduce_mulb1_ps12 ^ multm_reduce_mulb1_pc12;
  assign multm_reduce_vs13 = multm_reduce_mulb1_ps13 ^ multm_reduce_mulb1_pc13;
  assign multm_reduce_vs14 = multm_reduce_mulb1_ps14 ^ multm_reduce_mulb1_pc14;
  assign multm_reduce_vs15 = multm_reduce_mulb1_ps15 ^ multm_reduce_mulb1_pc15;
  assign multm_reduce_vs16 = multm_reduce_mulb1_ps16 ^ multm_reduce_mulb1_pc16;
  assign multm_reduce_vs17 = multm_reduce_mulb1_ps17 ^ multm_reduce_mulb1_pc17;
  assign multm_reduce_vs18 = multm_reduce_mulb1_ps18 ^ multm_reduce_mulb1_pc18;
  assign multm_reduce_vs19 = multm_reduce_mulb1_ps19 ^ multm_reduce_mulb1_pc19;
  assign multm_reduce_vs20 = multm_reduce_mulb1_ps20 ^ multm_reduce_mulb1_pc20;
  assign multm_reduce_vs21 = multm_reduce_mulb1_ps21 ^ multm_reduce_mulb1_pc21;
  assign multm_reduce_vs22 = multm_reduce_mulb1_ps22 ^ multm_reduce_mulb1_pc22;
  assign multm_reduce_vs23 = multm_reduce_mulb1_ps23 ^ multm_reduce_mulb1_pc23;
  assign multm_reduce_vs24 = multm_reduce_mulb1_ps24 ^ multm_reduce_mulb1_pc24;
  assign multm_reduce_vs25 = multm_reduce_mulb1_ps25 ^ multm_reduce_mulb1_pc25;
  assign multm_reduce_vs26 = multm_reduce_mulb1_ps26 ^ multm_reduce_mulb1_pc26;
  assign multm_reduce_vs27 = multm_reduce_mulb1_ps27 ^ multm_reduce_mulb1_pc27;
  assign multm_reduce_vs28 = multm_reduce_mulb1_ps28 ^ multm_reduce_mulb1_pc28;
  assign multm_reduce_vs29 = multm_reduce_mulb1_ps29 ^ multm_reduce_mulb1_pc29;
  assign multm_reduce_vs30 = multm_reduce_mulb1_ps30 ^ multm_reduce_mulb1_pc30;
  assign multm_reduce_vs31 = multm_reduce_mulb1_ps31 ^ multm_reduce_mulb1_pc31;
  assign multm_reduce_vs32 = multm_reduce_mulb1_ps32 ^ multm_reduce_mulb1_pc32;
  assign multm_reduce_vs33 = multm_reduce_mulb1_ps33 ^ multm_reduce_mulb1_pc33;
  assign multm_reduce_vs34 = multm_reduce_mulb1_ps34 ^ multm_reduce_mulb1_pc34;
  assign multm_reduce_vs35 = multm_reduce_mulb1_ps35 ^ multm_reduce_mulb1_pc35;
  assign multm_reduce_vs36 = multm_reduce_mulb1_ps36 ^ multm_reduce_mulb1_pc36;
  assign multm_reduce_vs37 = multm_reduce_mulb1_ps37 ^ multm_reduce_mulb1_pc37;
  assign multm_reduce_vs38 = multm_reduce_mulb1_ps38 ^ multm_reduce_mulb1_pc38;
  assign multm_reduce_vs39 = multm_reduce_mulb1_ps39 ^ multm_reduce_mulb1_pc39;
  assign multm_reduce_vs40 = multm_reduce_mulb1_ps40 ^ multm_reduce_mulb1_pc40;
  assign multm_reduce_vs41 = multm_reduce_mulb1_ps41 ^ multm_reduce_mulb1_pc41;
  assign multm_reduce_vs42 = multm_reduce_mulb1_ps42 ^ multm_reduce_mulb1_pc42;
  assign multm_reduce_vs43 = multm_reduce_mulb1_ps43 ^ multm_reduce_mulb1_pc43;
  assign multm_reduce_vs44 = multm_reduce_mulb1_ps44 ^ multm_reduce_mulb1_pc44;
  assign multm_reduce_vs45 = multm_reduce_mulb1_ps45 ^ multm_reduce_mulb1_pc45;
  assign multm_reduce_vs46 = multm_reduce_mulb1_ps46 ^ multm_reduce_mulb1_pc46;
  assign multm_reduce_vs47 = multm_reduce_mulb1_ps47 ^ multm_reduce_mulb1_pc47;
  assign multm_reduce_vs48 = multm_reduce_mulb1_ps48 ^ multm_reduce_mulb1_pc48;
  assign multm_reduce_vs49 = multm_reduce_mulb1_ps49 ^ multm_reduce_mulb1_pc49;
  assign multm_reduce_vs50 = multm_reduce_mulb1_ps50 ^ multm_reduce_mulb1_pc50;
  assign multm_reduce_vs51 = multm_reduce_mulb1_ps51 ^ multm_reduce_mulb1_pc51;
  assign multm_reduce_vs52 = multm_reduce_mulb1_ps52 ^ multm_reduce_mulb1_pc52;
  assign multm_reduce_vs53 = multm_reduce_mulb1_ps53 ^ multm_reduce_mulb1_pc53;
  assign multm_reduce_vs54 = multm_reduce_mulb1_ps54 ^ multm_reduce_mulb1_pc54;
  assign multm_reduce_vs55 = multm_reduce_mulb1_ps55 ^ multm_reduce_mulb1_pc55;
  assign multm_reduce_vs56 = multm_reduce_mulb1_ps56 ^ multm_reduce_mulb1_pc56;
  assign multm_reduce_vs57 = multm_reduce_mulb1_ps57 ^ multm_reduce_mulb1_pc57;
  assign multm_reduce_vs58 = multm_reduce_mulb1_ps58 ^ multm_reduce_mulb1_pc58;
  assign multm_reduce_vs59 = multm_reduce_mulb1_ps59 ^ multm_reduce_mulb1_pc59;
  assign multm_reduce_vs60 = multm_reduce_mulb1_ps60 ^ multm_reduce_mulb1_pc60;
  assign multm_reduce_vs61 = multm_reduce_mulb1_ps61 ^ multm_reduce_mulb1_pc61;
  assign multm_reduce_vs62 = multm_reduce_mulb1_ps62 ^ multm_reduce_mulb1_pc62;
  assign multm_reduce_vs63 = multm_reduce_mulb1_ps63 ^ multm_reduce_mulb1_pc63;
  assign multm_reduce_vs64 = multm_reduce_mulb1_ps64 ^ multm_reduce_mulb1_pc64;
  assign multm_reduce_vs65 = multm_reduce_mulb1_ps65 ^ multm_reduce_mulb1_pc65;
  assign multm_reduce_vs66 = multm_reduce_mulb1_ps66 ^ multm_reduce_mulb1_pc66;
  assign multm_reduce_vs67 = multm_reduce_mulb1_ps67 ^ multm_reduce_mulb1_pc67;
  assign multm_reduce_vs68 = multm_reduce_mulb1_ps68 ^ multm_reduce_mulb1_pc68;
  assign multm_reduce_vs69 = multm_reduce_mulb1_ps69 ^ multm_reduce_mulb1_pc69;
  assign multm_reduce_vs70 = multm_reduce_mulb1_ps70 ^ multm_reduce_mulb1_pc70;
  assign multm_reduce_vs71 = multm_reduce_mulb1_ps71 ^ multm_reduce_mulb1_pc71;
  assign multm_reduce_vs72 = multm_reduce_mulb1_ps72 ^ multm_reduce_mulb1_pc72;
  assign multm_reduce_vs73 = multm_reduce_mulb1_ps73 ^ multm_reduce_mulb1_pc73;
  assign multm_reduce_vs74 = multm_reduce_mulb1_ps74 ^ multm_reduce_mulb1_pc74;
  assign multm_reduce_vs75 = multm_reduce_mulb1_ps75 ^ multm_reduce_mulb1_pc75;
  assign multm_reduce_vs76 = multm_reduce_mulb1_ps76 ^ multm_reduce_mulb1_pc76;
  assign multm_reduce_vs77 = multm_reduce_mulb1_ps77 ^ multm_reduce_mulb1_pc77;
  assign multm_reduce_vs78 = multm_reduce_mulb1_ps78 ^ multm_reduce_mulb1_pc78;
  assign multm_reduce_vs79 = multm_reduce_mulb1_ps79 ^ multm_reduce_mulb1_pc79;
  assign multm_reduce_vs80 = multm_reduce_mulb1_ps80 ^ multm_reduce_mulb1_pc80;
  assign multm_reduce_vs81 = multm_reduce_mulb1_ps81 ^ multm_reduce_mulb1_pc81;
  assign multm_reduce_vs82 = multm_reduce_mulb1_ps82 ^ multm_reduce_mulb1_pc82;
  assign multm_reduce_vs83 = multm_reduce_mulb1_ps83 ^ multm_reduce_mulb1_pc83;
  assign multm_reduce_vs84 = multm_reduce_mulb1_ps84 ^ multm_reduce_mulb1_pc84;
  assign multm_reduce_vs85 = multm_reduce_mulb1_ps85 ^ multm_reduce_mulb1_pc85;
  assign multm_reduce_vs86 = multm_reduce_mulb1_ps86 ^ multm_reduce_mulb1_pc86;
  assign multm_reduce_vs87 = multm_reduce_mulb1_ps87 ^ multm_reduce_mulb1_pc87;
  assign multm_reduce_vs88 = multm_reduce_mulb1_ps88 ^ multm_reduce_mulb1_pc88;
  assign multm_reduce_vs89 = multm_reduce_mulb1_ps89 ^ multm_reduce_mulb1_pc89;
  assign multm_reduce_vs90 = multm_reduce_mulb1_ps90 ^ multm_reduce_mulb1_pc90;
  assign multm_reduce_vs91 = multm_reduce_mulb1_ps91 ^ multm_reduce_mulb1_pc91;
  assign multm_reduce_vs92 = multm_reduce_mulb1_ps92 ^ multm_reduce_mulb1_pc92;
  assign multm_reduce_vs93 = multm_reduce_mulb1_ps93 ^ multm_reduce_mulb1_pc93;
  assign multm_reduce_vs94 = multm_reduce_mulb1_ps94 ^ multm_reduce_mulb1_pc94;
  assign multm_reduce_vs95 = multm_reduce_mulb1_ps95 ^ multm_reduce_mulb1_pc95;
  assign multm_reduce_vs96 = multm_reduce_mulb1_ps96 ^ multm_reduce_mulb1_pc96;
  assign multm_reduce_vs97 = multm_reduce_mulb1_ps97 ^ multm_reduce_mulb1_pc97;
  assign multm_reduce_vs98 = multm_reduce_mulb1_ps98 ^ multm_reduce_mulb1_pc98;
  assign multm_reduce_vs99 = multm_reduce_mulb1_ps99 ^ multm_reduce_mulb1_pc99;
  assign multm_reduce_vs100 = multm_reduce_mulb1_ps100 ^ multm_reduce_mulb1_pc100;
  assign multm_reduce_vs101 = multm_reduce_mulb1_ps101 ^ multm_reduce_mulb1_pc101;
  assign multm_reduce_vs102 = multm_reduce_mulb1_ps102 ^ multm_reduce_mulb1_pc102;
  assign multm_reduce_vs103 = multm_reduce_mulb1_ps103 ^ multm_reduce_mulb1_pc103;
  assign multm_reduce_vs104 = multm_reduce_mulb1_ps104 ^ multm_reduce_mulb1_pc104;
  assign multm_reduce_vs105 = multm_reduce_mulb1_ps105 ^ multm_reduce_mulb1_pc105;
  assign multm_reduce_vs106 = multm_reduce_mulb1_ps106 ^ multm_reduce_mulb1_pc106;
  assign multm_reduce_vs107 = multm_reduce_mulb1_ps107 ^ multm_reduce_mulb1_pc107;
  assign multm_reduce_vs108 = multm_reduce_mulb1_ps108 ^ multm_reduce_mulb1_pc108;
  assign multm_reduce_vs109 = multm_reduce_mulb1_ps109 ^ multm_reduce_mulb1_pc109;
  assign multm_reduce_vs110 = multm_reduce_mulb1_ps110 ^ multm_reduce_mulb1_pc110;
  assign multm_reduce_vs111 = multm_reduce_mulb1_ps111 ^ multm_reduce_mulb1_pc111;
  assign multm_reduce_vs112 = multm_reduce_mulb1_ps112 ^ multm_reduce_mulb1_pc112;
  assign multm_reduce_vs113 = multm_reduce_mulb1_ps113 ^ multm_reduce_mulb1_pc113;
  assign multm_reduce_vs114 = multm_reduce_mulb1_ps114 ^ multm_reduce_mulb1_pc114;
  assign multm_reduce_vs115 = multm_reduce_mulb1_ps115 ^ multm_reduce_mulb1_pc115;
  assign multm_reduce_vs116 = multm_reduce_mulb1_ps116 ^ multm_reduce_mulb1_pc116;
  assign multm_reduce_vs117 = multm_reduce_mulb1_ps117 ^ multm_reduce_mulb1_pc117;
  assign multm_reduce_vs118 = multm_reduce_mulb1_ps118 ^ multm_reduce_mulb1_pc118;
  assign multm_reduce_vs119 = multm_reduce_mulb1_ps119 ^ multm_reduce_mulb1_pc119;
  assign multm_reduce_vs120 = multm_reduce_mulb1_ps120 ^ multm_reduce_mulb1_pc120;
  assign multm_reduce_vs121 = multm_reduce_mulb1_ps121 ^ multm_reduce_mulb1_pc121;
  assign multm_reduce_vs122 = multm_reduce_mulb1_ps122 ^ multm_reduce_mulb1_pc122;
  assign multm_reduce_vs123 = multm_reduce_mulb1_ps123 ^ multm_reduce_mulb1_pc123;
  assign multm_reduce_vs124 = multm_reduce_mulb1_ps124 ^ multm_reduce_mulb1_pc124;
  assign multm_reduce_vs125 = multm_reduce_mulb1_ps125 ^ multm_reduce_mulb1_pc125;
  assign multm_reduce_vs126 = multm_reduce_mulb1_ps126 ^ multm_reduce_mulb1_pc126;
  assign multm_reduce_vs127 = multm_reduce_mulb1_ps127 ^ multm_reduce_mulb1_pc127;
  assign multm_reduce_vs128 = multm_reduce_mulb1_ps128 ^ multm_reduce_mulb1_pc128;
  assign multm_reduce_vs129 = multm_reduce_mulb1_ps129 ^ multm_reduce_mulb1_pc129;
  assign multm_reduce_vs130 = multm_reduce_mulb1_ps130 ^ multm_reduce_mulb1_pc130;
  assign multm_reduce_vs131 = multm_reduce_mulb1_ps131 ^ multm_reduce_mulb1_pc131;
  assign multm_reduce_vs132 = multm_reduce_mulb1_ps132 ^ multm_reduce_mulb1_pc132;
  assign multm_reduce_vs133 = multm_reduce_mulb1_ps133 ^ multm_reduce_mulb1_pc133;
  assign multm_reduce_vs134 = multm_reduce_mulb1_ps134 ^ multm_reduce_mulb1_pc134;
  assign multm_reduce_vs135 = multm_reduce_mulb1_ps135 ^ multm_reduce_mulb1_pc135;
  assign multm_reduce_vs136 = multm_reduce_mulb1_ps136 ^ multm_reduce_mulb1_pc136;
  assign multm_reduce_vs137 = multm_reduce_mulb1_ps137 ^ multm_reduce_mulb1_pc137;
  assign multm_reduce_vs138 = multm_reduce_mulb1_ps138 ^ multm_reduce_mulb1_pc138;
  assign multm_reduce_vs139 = multm_reduce_mulb1_ps139 ^ multm_reduce_mulb1_pc139;
  assign multm_reduce_vs140 = multm_reduce_mulb1_ps140 ^ multm_reduce_mulb1_pc140;
  assign multm_reduce_vs141 = multm_reduce_mulb1_ps141 ^ multm_reduce_mulb1_pc141;
  assign multm_reduce_vs142 = multm_reduce_mulb1_ps142 ^ multm_reduce_mulb1_pc142;
  assign multm_reduce_vs143 = multm_reduce_mulb1_ps143 ^ multm_reduce_mulb1_pc143;
  assign multm_reduce_vs144 = multm_reduce_mulb1_ps144 ^ multm_reduce_mulb1_pc144;
  assign multm_reduce_vs145 = multm_reduce_mulb1_ps145 ^ multm_reduce_mulb1_pc145;
  assign multm_reduce_vs146 = multm_reduce_mulb1_ps146 ^ multm_reduce_mulb1_pc146;
  assign multm_reduce_vs147 = multm_reduce_mulb1_ps147 ^ multm_reduce_mulb1_pc147;
  assign multm_reduce_vs148 = multm_reduce_mulb1_ps148 ^ multm_reduce_mulb1_pc148;
  assign multm_reduce_vs149 = multm_reduce_mulb1_ps149 ^ multm_reduce_mulb1_pc149;
  assign multm_reduce_vs150 = multm_reduce_mulb1_ps150 ^ multm_reduce_mulb1_pc150;
  assign multm_reduce_vs151 = multm_reduce_mulb1_ps151 ^ multm_reduce_mulb1_pc151;
  assign multm_reduce_vs152 = multm_reduce_mulb1_ps152 ^ multm_reduce_mulb1_pc152;
  assign multm_reduce_vs153 = multm_reduce_mulb1_ps153 ^ multm_reduce_mulb1_pc153;
  assign multm_reduce_vs154 = multm_reduce_mulb1_ps154 ^ multm_reduce_mulb1_pc154;
  assign multm_reduce_vs155 = multm_reduce_mulb1_ps155 ^ multm_reduce_mulb1_pc155;
  assign multm_reduce_vs156 = multm_reduce_mulb1_ps156 ^ multm_reduce_mulb1_pc156;
  assign multm_reduce_vs157 = multm_reduce_mulb1_ps157 ^ multm_reduce_mulb1_pc157;
  assign multm_reduce_vs158 = multm_reduce_mulb1_ps158 ^ multm_reduce_mulb1_pc158;
  assign multm_reduce_vs159 = multm_reduce_mulb1_ps159 ^ multm_reduce_mulb1_pc159;
  assign multm_reduce_vs160 = multm_reduce_mulb1_ps160 ^ multm_reduce_mulb1_pc160;
  assign multm_reduce_vs161 = multm_reduce_mulb1_ps161 ^ multm_reduce_mulb1_pc161;
  assign multm_reduce_vs162 = multm_reduce_mulb1_ps162 ^ multm_reduce_mulb1_pc162;
  assign multm_reduce_vs163 = multm_reduce_mulb1_ps163 ^ multm_reduce_mulb1_pc163;
  assign multm_reduce_vs164 = multm_reduce_mulb1_ps164 ^ multm_reduce_mulb1_pc164;
  assign multm_reduce_vs165 = multm_reduce_mulb1_ps165 ^ multm_reduce_mulb1_pc165;
  assign multm_reduce_vs166 = multm_reduce_mulb1_ps166 ^ multm_reduce_mulb1_pc166;
  assign multm_reduce_vs167 = multm_reduce_mulb1_ps167 ^ multm_reduce_mulb1_pc167;
  assign multm_reduce_vs168 = multm_reduce_mulb1_ps168 ^ multm_reduce_mulb1_pc168;
  assign multm_reduce_vs169 = multm_reduce_mulb1_ps169 ^ multm_reduce_mulb1_pc169;
  assign multm_reduce_vs170 = multm_reduce_mulb1_ps170 ^ multm_reduce_mulb1_pc170;
  assign multm_reduce_vs171 = multm_reduce_mulb1_ps171 ^ multm_reduce_mulb1_pc171;
  assign multm_reduce_vs172 = multm_reduce_mulb1_ps172 ^ multm_reduce_mulb1_pc172;
  assign multm_reduce_vs173 = multm_reduce_mulb1_ps173 ^ multm_reduce_mulb1_pc173;
  assign multm_reduce_vs174 = multm_reduce_mulb1_ps174 ^ multm_reduce_mulb1_pc174;
  assign multm_reduce_vs175 = multm_reduce_mulb1_ps175 ^ multm_reduce_mulb1_pc175;
  assign multm_reduce_vs176 = multm_reduce_mulb1_ps176 ^ multm_reduce_mulb1_pc176;
  assign multm_reduce_vs177 = multm_reduce_mulb1_ps177 ^ multm_reduce_mulb1_pc177;
  assign multm_reduce_vs178 = multm_reduce_mulb1_ps178 ^ multm_reduce_mulb1_pc178;
  assign multm_reduce_vs179 = multm_reduce_mulb1_ps179 ^ multm_reduce_mulb1_pc179;
  assign multm_reduce_vs180 = multm_reduce_mulb1_ps180 ^ multm_reduce_mulb1_pc180;
  assign multm_reduce_vs181 = multm_reduce_mulb1_ps181 ^ multm_reduce_mulb1_pc181;
  assign multm_reduce_vs182 = multm_reduce_mulb1_add3_xor3_wx ^ multm_reduce_mulb1_pc182;
  assign multm_reduce_vt = multm_reduce_vb | multm_reduce_sticky_q;
  assign nor2_zn = sad | sbd;
  assign pcq0 = sbd ? xc[0] : qc0;
  assign pcq1 = sbd ? xc[1] : qc1;
  assign pcq2 = sbd ? xc[2] : qc2;
  assign pcq3 = sbd ? xc[3] : qc3;
  assign pcq4 = sbd ? xc[4] : qc4;
  assign pcq5 = sbd ? xc[5] : qc5;
  assign pcq6 = sbd ? xc[6] : qc6;
  assign pcq7 = sbd ? xc[7] : qc7;
  assign pcq8 = sbd ? xc[8] : qc8;
  assign pcq9 = sbd ? xc[9] : qc9;
  assign pcq10 = sbd ? xc[10] : qc10;
  assign pcq11 = sbd ? xc[11] : qc11;
  assign pcq12 = sbd ? xc[12] : qc12;
  assign pcq13 = sbd ? xc[13] : qc13;
  assign pcq14 = sbd ? xc[14] : qc14;
  assign pcq15 = sbd ? xc[15] : qc15;
  assign pcq16 = sbd ? xc[16] : qc16;
  assign pcq17 = sbd ? xc[17] : qc17;
  assign pcq18 = sbd ? xc[18] : qc18;
  assign pcq19 = sbd ? xc[19] : qc19;
  assign pcq20 = sbd ? xc[20] : qc20;
  assign pcq21 = sbd ? xc[21] : qc21;
  assign pcq22 = sbd ? xc[22] : qc22;
  assign pcq23 = sbd ? xc[23] : qc23;
  assign pcq24 = sbd ? xc[24] : qc24;
  assign pcq25 = sbd ? xc[25] : qc25;
  assign pcq26 = sbd ? xc[26] : qc26;
  assign pcq27 = sbd ? xc[27] : qc27;
  assign pcq28 = sbd ? xc[28] : qc28;
  assign pcq29 = sbd ? xc[29] : qc29;
  assign pcq30 = sbd ? xc[30] : qc30;
  assign pcq31 = sbd ? xc[31] : qc31;
  assign pcq32 = sbd ? xc[32] : qc32;
  assign pcq33 = sbd ? xc[33] : qc33;
  assign pcq34 = sbd ? xc[34] : qc34;
  assign pcq35 = sbd ? xc[35] : qc35;
  assign pcq36 = sbd ? xc[36] : qc36;
  assign pcq37 = sbd ? xc[37] : qc37;
  assign pcq38 = sbd ? xc[38] : qc38;
  assign pcq39 = sbd ? xc[39] : qc39;
  assign pcq40 = sbd ? xc[40] : qc40;
  assign pcq41 = sbd ? xc[41] : qc41;
  assign pcq42 = sbd ? xc[42] : qc42;
  assign pcq43 = sbd ? xc[43] : qc43;
  assign pcq44 = sbd ? xc[44] : qc44;
  assign pcq45 = sbd ? xc[45] : qc45;
  assign pcq46 = sbd ? xc[46] : qc46;
  assign pcq47 = sbd ? xc[47] : qc47;
  assign pcq48 = sbd ? xc[48] : qc48;
  assign pcq49 = sbd ? xc[49] : qc49;
  assign pcq50 = sbd ? xc[50] : qc50;
  assign pcq51 = sbd ? xc[51] : qc51;
  assign pcq52 = sbd ? xc[52] : qc52;
  assign pcq53 = sbd ? xc[53] : qc53;
  assign pcq54 = sbd ? xc[54] : qc54;
  assign pcq55 = sbd ? xc[55] : qc55;
  assign pcq56 = sbd ? xc[56] : qc56;
  assign pcq57 = sbd ? xc[57] : qc57;
  assign pcq58 = sbd ? xc[58] : qc58;
  assign pcq59 = sbd ? xc[59] : qc59;
  assign pcq60 = sbd ? xc[60] : qc60;
  assign pcq61 = sbd ? xc[61] : qc61;
  assign pcq62 = sbd ? xc[62] : qc62;
  assign pcq63 = sbd ? xc[63] : qc63;
  assign pcq64 = sbd ? xc[64] : qc64;
  assign pcq65 = sbd ? xc[65] : qc65;
  assign pcq66 = sbd ? xc[66] : qc66;
  assign pcq67 = sbd ? xc[67] : qc67;
  assign pcq68 = sbd ? xc[68] : qc68;
  assign pcq69 = sbd ? xc[69] : qc69;
  assign pcq70 = sbd ? xc[70] : qc70;
  assign pcq71 = sbd ? xc[71] : qc71;
  assign pcq72 = sbd ? xc[72] : qc72;
  assign pcq73 = sbd ? xc[73] : qc73;
  assign pcq74 = sbd ? xc[74] : qc74;
  assign pcq75 = sbd ? xc[75] : qc75;
  assign pcq76 = sbd ? xc[76] : qc76;
  assign pcq77 = sbd ? xc[77] : qc77;
  assign pcq78 = sbd ? xc[78] : qc78;
  assign pcq79 = sbd ? xc[79] : qc79;
  assign pcq80 = sbd ? xc[80] : qc80;
  assign pcq81 = sbd ? xc[81] : qc81;
  assign pcq82 = sbd ? xc[82] : qc82;
  assign pcq83 = sbd ? xc[83] : qc83;
  assign pcq84 = sbd ? xc[84] : qc84;
  assign pcq85 = sbd ? xc[85] : qc85;
  assign pcq86 = sbd ? xc[86] : qc86;
  assign pcq87 = sbd ? xc[87] : qc87;
  assign pcq88 = sbd ? xc[88] : qc88;
  assign pcq89 = sbd ? xc[89] : qc89;
  assign pcq90 = sbd ? xc[90] : qc90;
  assign pcq91 = sbd ? xc[91] : qc91;
  assign pcq92 = sbd ? xc[92] : qc92;
  assign pcq93 = sbd ? xc[93] : qc93;
  assign pcq94 = sbd ? xc[94] : qc94;
  assign pcq95 = sbd ? xc[95] : qc95;
  assign pcq96 = sbd ? xc[96] : qc96;
  assign pcq97 = sbd ? xc[97] : qc97;
  assign pcq98 = sbd ? xc[98] : qc98;
  assign pcq99 = sbd ? xc[99] : qc99;
  assign pcq100 = sbd ? xc[100] : qc100;
  assign pcq101 = sbd ? xc[101] : qc101;
  assign pcq102 = sbd ? xc[102] : qc102;
  assign pcq103 = sbd ? xc[103] : qc103;
  assign pcq104 = sbd ? xc[104] : qc104;
  assign pcq105 = sbd ? xc[105] : qc105;
  assign pcq106 = sbd ? xc[106] : qc106;
  assign pcq107 = sbd ? xc[107] : qc107;
  assign pcq108 = sbd ? xc[108] : qc108;
  assign pcq109 = sbd ? xc[109] : qc109;
  assign pcq110 = sbd ? xc[110] : qc110;
  assign pcq111 = sbd ? xc[111] : qc111;
  assign pcq112 = sbd ? xc[112] : qc112;
  assign pcq113 = sbd ? xc[113] : qc113;
  assign pcq114 = sbd ? xc[114] : qc114;
  assign pcq115 = sbd ? xc[115] : qc115;
  assign pcq116 = sbd ? xc[116] : qc116;
  assign pcq117 = sbd ? xc[117] : qc117;
  assign pcq118 = sbd ? xc[118] : qc118;
  assign pcq119 = sbd ? xc[119] : qc119;
  assign pcq120 = sbd ? xc[120] : qc120;
  assign pcq121 = sbd ? xc[121] : qc121;
  assign pcq122 = sbd ? xc[122] : qc122;
  assign pcq123 = sbd ? xc[123] : qc123;
  assign pcq124 = sbd ? xc[124] : qc124;
  assign pcq125 = sbd ? xc[125] : qc125;
  assign pcq126 = sbd ? xc[126] : qc126;
  assign pcq127 = sbd ? xc[127] : qc127;
  assign pcq128 = sbd ? xc[128] : qc128;
  assign pcq129 = sbd ? xc[129] : qc129;
  assign pcq130 = sbd ? xc[130] : qc130;
  assign pcq131 = sbd ? xc[131] : qc131;
  assign pcq132 = sbd ? xc[132] : qc132;
  assign pcq133 = sbd ? xc[133] : qc133;
  assign pcq134 = sbd ? xc[134] : qc134;
  assign pcq135 = sbd ? xc[135] : qc135;
  assign pcq136 = sbd ? xc[136] : qc136;
  assign pcq137 = sbd ? xc[137] : qc137;
  assign pcq138 = sbd ? xc[138] : qc138;
  assign pcq139 = sbd ? xc[139] : qc139;
  assign pcq140 = sbd ? xc[140] : qc140;
  assign pcq141 = sbd ? xc[141] : qc141;
  assign pcq142 = sbd ? xc[142] : qc142;
  assign pcq143 = sbd ? xc[143] : qc143;
  assign pcq144 = sbd ? xc[144] : qc144;
  assign pcq145 = sbd ? xc[145] : qc145;
  assign pcq146 = sbd ? xc[146] : qc146;
  assign pcq147 = sbd ? xc[147] : qc147;
  assign pcq148 = sbd ? xc[148] : qc148;
  assign pcq149 = sbd ? xc[149] : qc149;
  assign pcq150 = sbd ? xc[150] : qc150;
  assign pcq151 = sbd ? xc[151] : qc151;
  assign pcq152 = sbd ? xc[152] : qc152;
  assign pcq153 = sbd ? xc[153] : qc153;
  assign pcq154 = sbd ? xc[154] : qc154;
  assign pcq155 = sbd ? xc[155] : qc155;
  assign pcq156 = sbd ? xc[156] : qc156;
  assign pcq157 = sbd ? xc[157] : qc157;
  assign pcq158 = sbd ? xc[158] : qc158;
  assign pcq159 = sbd ? xc[159] : qc159;
  assign pcq160 = sbd ? xc[160] : qc160;
  assign pcq161 = sbd ? xc[161] : qc161;
  assign pcq162 = sbd ? xc[162] : qc162;
  assign pcq163 = sbd ? xc[163] : qc163;
  assign pcq164 = sbd ? xc[164] : qc164;
  assign pcq165 = sbd ? xc[165] : qc165;
  assign pcq166 = sbd ? xc[166] : qc166;
  assign pcq167 = sbd ? xc[167] : qc167;
  assign pcq168 = sbd ? xc[168] : qc168;
  assign pcq169 = sbd ? xc[169] : qc169;
  assign pcq170 = sbd ? xc[170] : qc170;
  assign pcq171 = sbd ? xc[171] : qc171;
  assign pcq172 = sbd ? xc[172] : qc172;
  assign pcq173 = sbd ? xc[173] : qc173;
  assign pcq174 = sbd ? xc[174] : qc174;
  assign pcq175 = sbd ? xc[175] : qc175;
  assign pcq176 = sbd ? xc[176] : qc176;
  assign pcq177 = sbd ? xc[177] : qc177;
  assign pcq178 = sbd ? xc[178] : qc178;
  assign pcq179 = sbd ? xc[179] : qc179;
  assign pcq180 = sbd ? xc[180] : qc180;
  assign pcq181 = sbd ? xc[181] : qc181;
  assign pcq182 = sbd ? xc[182] : qc182;
  assign pcq183 = sbd ? xc[183] : qc183;
  assign pcr0 = sad ? pcq0 : yc0_o;
  assign pcr1 = sad ? pcq1 : yc1_o;
  assign pcr2 = sad ? pcq2 : yc2_o;
  assign pcr3 = sad ? pcq3 : yc3_o;
  assign pcr4 = sad ? pcq4 : yc4_o;
  assign pcr5 = sad ? pcq5 : yc5_o;
  assign pcr6 = sad ? pcq6 : yc6_o;
  assign pcr7 = sad ? pcq7 : yc7_o;
  assign pcr8 = sad ? pcq8 : yc8_o;
  assign pcr9 = sad ? pcq9 : yc9_o;
  assign pcr10 = sad ? pcq10 : yc10_o;
  assign pcr11 = sad ? pcq11 : yc11_o;
  assign pcr12 = sad ? pcq12 : yc12_o;
  assign pcr13 = sad ? pcq13 : yc13_o;
  assign pcr14 = sad ? pcq14 : yc14_o;
  assign pcr15 = sad ? pcq15 : yc15_o;
  assign pcr16 = sad ? pcq16 : yc16_o;
  assign pcr17 = sad ? pcq17 : yc17_o;
  assign pcr18 = sad ? pcq18 : yc18_o;
  assign pcr19 = sad ? pcq19 : yc19_o;
  assign pcr20 = sad ? pcq20 : yc20_o;
  assign pcr21 = sad ? pcq21 : yc21_o;
  assign pcr22 = sad ? pcq22 : yc22_o;
  assign pcr23 = sad ? pcq23 : yc23_o;
  assign pcr24 = sad ? pcq24 : yc24_o;
  assign pcr25 = sad ? pcq25 : yc25_o;
  assign pcr26 = sad ? pcq26 : yc26_o;
  assign pcr27 = sad ? pcq27 : yc27_o;
  assign pcr28 = sad ? pcq28 : yc28_o;
  assign pcr29 = sad ? pcq29 : yc29_o;
  assign pcr30 = sad ? pcq30 : yc30_o;
  assign pcr31 = sad ? pcq31 : yc31_o;
  assign pcr32 = sad ? pcq32 : yc32_o;
  assign pcr33 = sad ? pcq33 : yc33_o;
  assign pcr34 = sad ? pcq34 : yc34_o;
  assign pcr35 = sad ? pcq35 : yc35_o;
  assign pcr36 = sad ? pcq36 : yc36_o;
  assign pcr37 = sad ? pcq37 : yc37_o;
  assign pcr38 = sad ? pcq38 : yc38_o;
  assign pcr39 = sad ? pcq39 : yc39_o;
  assign pcr40 = sad ? pcq40 : yc40_o;
  assign pcr41 = sad ? pcq41 : yc41_o;
  assign pcr42 = sad ? pcq42 : yc42_o;
  assign pcr43 = sad ? pcq43 : yc43_o;
  assign pcr44 = sad ? pcq44 : yc44_o;
  assign pcr45 = sad ? pcq45 : yc45_o;
  assign pcr46 = sad ? pcq46 : yc46_o;
  assign pcr47 = sad ? pcq47 : yc47_o;
  assign pcr48 = sad ? pcq48 : yc48_o;
  assign pcr49 = sad ? pcq49 : yc49_o;
  assign pcr50 = sad ? pcq50 : yc50_o;
  assign pcr51 = sad ? pcq51 : yc51_o;
  assign pcr52 = sad ? pcq52 : yc52_o;
  assign pcr53 = sad ? pcq53 : yc53_o;
  assign pcr54 = sad ? pcq54 : yc54_o;
  assign pcr55 = sad ? pcq55 : yc55_o;
  assign pcr56 = sad ? pcq56 : yc56_o;
  assign pcr57 = sad ? pcq57 : yc57_o;
  assign pcr58 = sad ? pcq58 : yc58_o;
  assign pcr59 = sad ? pcq59 : yc59_o;
  assign pcr60 = sad ? pcq60 : yc60_o;
  assign pcr61 = sad ? pcq61 : yc61_o;
  assign pcr62 = sad ? pcq62 : yc62_o;
  assign pcr63 = sad ? pcq63 : yc63_o;
  assign pcr64 = sad ? pcq64 : yc64_o;
  assign pcr65 = sad ? pcq65 : yc65_o;
  assign pcr66 = sad ? pcq66 : yc66_o;
  assign pcr67 = sad ? pcq67 : yc67_o;
  assign pcr68 = sad ? pcq68 : yc68_o;
  assign pcr69 = sad ? pcq69 : yc69_o;
  assign pcr70 = sad ? pcq70 : yc70_o;
  assign pcr71 = sad ? pcq71 : yc71_o;
  assign pcr72 = sad ? pcq72 : yc72_o;
  assign pcr73 = sad ? pcq73 : yc73_o;
  assign pcr74 = sad ? pcq74 : yc74_o;
  assign pcr75 = sad ? pcq75 : yc75_o;
  assign pcr76 = sad ? pcq76 : yc76_o;
  assign pcr77 = sad ? pcq77 : yc77_o;
  assign pcr78 = sad ? pcq78 : yc78_o;
  assign pcr79 = sad ? pcq79 : yc79_o;
  assign pcr80 = sad ? pcq80 : yc80_o;
  assign pcr81 = sad ? pcq81 : yc81_o;
  assign pcr82 = sad ? pcq82 : yc82_o;
  assign pcr83 = sad ? pcq83 : yc83_o;
  assign pcr84 = sad ? pcq84 : yc84_o;
  assign pcr85 = sad ? pcq85 : yc85_o;
  assign pcr86 = sad ? pcq86 : yc86_o;
  assign pcr87 = sad ? pcq87 : yc87_o;
  assign pcr88 = sad ? pcq88 : yc88_o;
  assign pcr89 = sad ? pcq89 : yc89_o;
  assign pcr90 = sad ? pcq90 : yc90_o;
  assign pcr91 = sad ? pcq91 : yc91_o;
  assign pcr92 = sad ? pcq92 : yc92_o;
  assign pcr93 = sad ? pcq93 : yc93_o;
  assign pcr94 = sad ? pcq94 : yc94_o;
  assign pcr95 = sad ? pcq95 : yc95_o;
  assign pcr96 = sad ? pcq96 : yc96_o;
  assign pcr97 = sad ? pcq97 : yc97_o;
  assign pcr98 = sad ? pcq98 : yc98_o;
  assign pcr99 = sad ? pcq99 : yc99_o;
  assign pcr100 = sad ? pcq100 : yc100_o;
  assign pcr101 = sad ? pcq101 : yc101_o;
  assign pcr102 = sad ? pcq102 : yc102_o;
  assign pcr103 = sad ? pcq103 : yc103_o;
  assign pcr104 = sad ? pcq104 : yc104_o;
  assign pcr105 = sad ? pcq105 : yc105_o;
  assign pcr106 = sad ? pcq106 : yc106_o;
  assign pcr107 = sad ? pcq107 : yc107_o;
  assign pcr108 = sad ? pcq108 : yc108_o;
  assign pcr109 = sad ? pcq109 : yc109_o;
  assign pcr110 = sad ? pcq110 : yc110_o;
  assign pcr111 = sad ? pcq111 : yc111_o;
  assign pcr112 = sad ? pcq112 : yc112_o;
  assign pcr113 = sad ? pcq113 : yc113_o;
  assign pcr114 = sad ? pcq114 : yc114_o;
  assign pcr115 = sad ? pcq115 : yc115_o;
  assign pcr116 = sad ? pcq116 : yc116_o;
  assign pcr117 = sad ? pcq117 : yc117_o;
  assign pcr118 = sad ? pcq118 : yc118_o;
  assign pcr119 = sad ? pcq119 : yc119_o;
  assign pcr120 = sad ? pcq120 : yc120_o;
  assign pcr121 = sad ? pcq121 : yc121_o;
  assign pcr122 = sad ? pcq122 : yc122_o;
  assign pcr123 = sad ? pcq123 : yc123_o;
  assign pcr124 = sad ? pcq124 : yc124_o;
  assign pcr125 = sad ? pcq125 : yc125_o;
  assign pcr126 = sad ? pcq126 : yc126_o;
  assign pcr127 = sad ? pcq127 : yc127_o;
  assign pcr128 = sad ? pcq128 : yc128_o;
  assign pcr129 = sad ? pcq129 : yc129_o;
  assign pcr130 = sad ? pcq130 : yc130_o;
  assign pcr131 = sad ? pcq131 : yc131_o;
  assign pcr132 = sad ? pcq132 : yc132_o;
  assign pcr133 = sad ? pcq133 : yc133_o;
  assign pcr134 = sad ? pcq134 : yc134_o;
  assign pcr135 = sad ? pcq135 : yc135_o;
  assign pcr136 = sad ? pcq136 : yc136_o;
  assign pcr137 = sad ? pcq137 : yc137_o;
  assign pcr138 = sad ? pcq138 : yc138_o;
  assign pcr139 = sad ? pcq139 : yc139_o;
  assign pcr140 = sad ? pcq140 : yc140_o;
  assign pcr141 = sad ? pcq141 : yc141_o;
  assign pcr142 = sad ? pcq142 : yc142_o;
  assign pcr143 = sad ? pcq143 : yc143_o;
  assign pcr144 = sad ? pcq144 : yc144_o;
  assign pcr145 = sad ? pcq145 : yc145_o;
  assign pcr146 = sad ? pcq146 : yc146_o;
  assign pcr147 = sad ? pcq147 : yc147_o;
  assign pcr148 = sad ? pcq148 : yc148_o;
  assign pcr149 = sad ? pcq149 : yc149_o;
  assign pcr150 = sad ? pcq150 : yc150_o;
  assign pcr151 = sad ? pcq151 : yc151_o;
  assign pcr152 = sad ? pcq152 : yc152_o;
  assign pcr153 = sad ? pcq153 : yc153_o;
  assign pcr154 = sad ? pcq154 : yc154_o;
  assign pcr155 = sad ? pcq155 : yc155_o;
  assign pcr156 = sad ? pcq156 : yc156_o;
  assign pcr157 = sad ? pcq157 : yc157_o;
  assign pcr158 = sad ? pcq158 : yc158_o;
  assign pcr159 = sad ? pcq159 : yc159_o;
  assign pcr160 = sad ? pcq160 : yc160_o;
  assign pcr161 = sad ? pcq161 : yc161_o;
  assign pcr162 = sad ? pcq162 : yc162_o;
  assign pcr163 = sad ? pcq163 : yc163_o;
  assign pcr164 = sad ? pcq164 : yc164_o;
  assign pcr165 = sad ? pcq165 : yc165_o;
  assign pcr166 = sad ? pcq166 : yc166_o;
  assign pcr167 = sad ? pcq167 : yc167_o;
  assign pcr168 = sad ? pcq168 : yc168_o;
  assign pcr169 = sad ? pcq169 : yc169_o;
  assign pcr170 = sad ? pcq170 : yc170_o;
  assign pcr171 = sad ? pcq171 : yc171_o;
  assign pcr172 = sad ? pcq172 : yc172_o;
  assign pcr173 = sad ? pcq173 : yc173_o;
  assign pcr174 = sad ? pcq174 : yc174_o;
  assign pcr175 = sad ? pcq175 : yc175_o;
  assign pcr176 = sad ? pcq176 : yc176_o;
  assign pcr177 = sad ? pcq177 : yc177_o;
  assign pcr178 = sad ? pcq178 : yc178_o;
  assign pcr179 = sad ? pcq179 : yc179_o;
  assign pcr180 = sad ? pcq180 : yc180_o;
  assign pcr181 = sad ? pcq181 : yc181_o;
  assign pcr182 = sad ? pcq182 : yc182_o;
  assign pcr183 = sad ? pcq183 : yc183_o;
  assign psq0 = sbd ? xs[0] : qs0;
  assign psq1 = sbd ? xs[1] : qs1;
  assign psq2 = sbd ? xs[2] : qs2;
  assign psq3 = sbd ? xs[3] : qs3;
  assign psq4 = sbd ? xs[4] : qs4;
  assign psq5 = sbd ? xs[5] : qs5;
  assign psq6 = sbd ? xs[6] : qs6;
  assign psq7 = sbd ? xs[7] : qs7;
  assign psq8 = sbd ? xs[8] : qs8;
  assign psq9 = sbd ? xs[9] : qs9;
  assign psq10 = sbd ? xs[10] : qs10;
  assign psq11 = sbd ? xs[11] : qs11;
  assign psq12 = sbd ? xs[12] : qs12;
  assign psq13 = sbd ? xs[13] : qs13;
  assign psq14 = sbd ? xs[14] : qs14;
  assign psq15 = sbd ? xs[15] : qs15;
  assign psq16 = sbd ? xs[16] : qs16;
  assign psq17 = sbd ? xs[17] : qs17;
  assign psq18 = sbd ? xs[18] : qs18;
  assign psq19 = sbd ? xs[19] : qs19;
  assign psq20 = sbd ? xs[20] : qs20;
  assign psq21 = sbd ? xs[21] : qs21;
  assign psq22 = sbd ? xs[22] : qs22;
  assign psq23 = sbd ? xs[23] : qs23;
  assign psq24 = sbd ? xs[24] : qs24;
  assign psq25 = sbd ? xs[25] : qs25;
  assign psq26 = sbd ? xs[26] : qs26;
  assign psq27 = sbd ? xs[27] : qs27;
  assign psq28 = sbd ? xs[28] : qs28;
  assign psq29 = sbd ? xs[29] : qs29;
  assign psq30 = sbd ? xs[30] : qs30;
  assign psq31 = sbd ? xs[31] : qs31;
  assign psq32 = sbd ? xs[32] : qs32;
  assign psq33 = sbd ? xs[33] : qs33;
  assign psq34 = sbd ? xs[34] : qs34;
  assign psq35 = sbd ? xs[35] : qs35;
  assign psq36 = sbd ? xs[36] : qs36;
  assign psq37 = sbd ? xs[37] : qs37;
  assign psq38 = sbd ? xs[38] : qs38;
  assign psq39 = sbd ? xs[39] : qs39;
  assign psq40 = sbd ? xs[40] : qs40;
  assign psq41 = sbd ? xs[41] : qs41;
  assign psq42 = sbd ? xs[42] : qs42;
  assign psq43 = sbd ? xs[43] : qs43;
  assign psq44 = sbd ? xs[44] : qs44;
  assign psq45 = sbd ? xs[45] : qs45;
  assign psq46 = sbd ? xs[46] : qs46;
  assign psq47 = sbd ? xs[47] : qs47;
  assign psq48 = sbd ? xs[48] : qs48;
  assign psq49 = sbd ? xs[49] : qs49;
  assign psq50 = sbd ? xs[50] : qs50;
  assign psq51 = sbd ? xs[51] : qs51;
  assign psq52 = sbd ? xs[52] : qs52;
  assign psq53 = sbd ? xs[53] : qs53;
  assign psq54 = sbd ? xs[54] : qs54;
  assign psq55 = sbd ? xs[55] : qs55;
  assign psq56 = sbd ? xs[56] : qs56;
  assign psq57 = sbd ? xs[57] : qs57;
  assign psq58 = sbd ? xs[58] : qs58;
  assign psq59 = sbd ? xs[59] : qs59;
  assign psq60 = sbd ? xs[60] : qs60;
  assign psq61 = sbd ? xs[61] : qs61;
  assign psq62 = sbd ? xs[62] : qs62;
  assign psq63 = sbd ? xs[63] : qs63;
  assign psq64 = sbd ? xs[64] : qs64;
  assign psq65 = sbd ? xs[65] : qs65;
  assign psq66 = sbd ? xs[66] : qs66;
  assign psq67 = sbd ? xs[67] : qs67;
  assign psq68 = sbd ? xs[68] : qs68;
  assign psq69 = sbd ? xs[69] : qs69;
  assign psq70 = sbd ? xs[70] : qs70;
  assign psq71 = sbd ? xs[71] : qs71;
  assign psq72 = sbd ? xs[72] : qs72;
  assign psq73 = sbd ? xs[73] : qs73;
  assign psq74 = sbd ? xs[74] : qs74;
  assign psq75 = sbd ? xs[75] : qs75;
  assign psq76 = sbd ? xs[76] : qs76;
  assign psq77 = sbd ? xs[77] : qs77;
  assign psq78 = sbd ? xs[78] : qs78;
  assign psq79 = sbd ? xs[79] : qs79;
  assign psq80 = sbd ? xs[80] : qs80;
  assign psq81 = sbd ? xs[81] : qs81;
  assign psq82 = sbd ? xs[82] : qs82;
  assign psq83 = sbd ? xs[83] : qs83;
  assign psq84 = sbd ? xs[84] : qs84;
  assign psq85 = sbd ? xs[85] : qs85;
  assign psq86 = sbd ? xs[86] : qs86;
  assign psq87 = sbd ? xs[87] : qs87;
  assign psq88 = sbd ? xs[88] : qs88;
  assign psq89 = sbd ? xs[89] : qs89;
  assign psq90 = sbd ? xs[90] : qs90;
  assign psq91 = sbd ? xs[91] : qs91;
  assign psq92 = sbd ? xs[92] : qs92;
  assign psq93 = sbd ? xs[93] : qs93;
  assign psq94 = sbd ? xs[94] : qs94;
  assign psq95 = sbd ? xs[95] : qs95;
  assign psq96 = sbd ? xs[96] : qs96;
  assign psq97 = sbd ? xs[97] : qs97;
  assign psq98 = sbd ? xs[98] : qs98;
  assign psq99 = sbd ? xs[99] : qs99;
  assign psq100 = sbd ? xs[100] : qs100;
  assign psq101 = sbd ? xs[101] : qs101;
  assign psq102 = sbd ? xs[102] : qs102;
  assign psq103 = sbd ? xs[103] : qs103;
  assign psq104 = sbd ? xs[104] : qs104;
  assign psq105 = sbd ? xs[105] : qs105;
  assign psq106 = sbd ? xs[106] : qs106;
  assign psq107 = sbd ? xs[107] : qs107;
  assign psq108 = sbd ? xs[108] : qs108;
  assign psq109 = sbd ? xs[109] : qs109;
  assign psq110 = sbd ? xs[110] : qs110;
  assign psq111 = sbd ? xs[111] : qs111;
  assign psq112 = sbd ? xs[112] : qs112;
  assign psq113 = sbd ? xs[113] : qs113;
  assign psq114 = sbd ? xs[114] : qs114;
  assign psq115 = sbd ? xs[115] : qs115;
  assign psq116 = sbd ? xs[116] : qs116;
  assign psq117 = sbd ? xs[117] : qs117;
  assign psq118 = sbd ? xs[118] : qs118;
  assign psq119 = sbd ? xs[119] : qs119;
  assign psq120 = sbd ? xs[120] : qs120;
  assign psq121 = sbd ? xs[121] : qs121;
  assign psq122 = sbd ? xs[122] : qs122;
  assign psq123 = sbd ? xs[123] : qs123;
  assign psq124 = sbd ? xs[124] : qs124;
  assign psq125 = sbd ? xs[125] : qs125;
  assign psq126 = sbd ? xs[126] : qs126;
  assign psq127 = sbd ? xs[127] : qs127;
  assign psq128 = sbd ? xs[128] : qs128;
  assign psq129 = sbd ? xs[129] : qs129;
  assign psq130 = sbd ? xs[130] : qs130;
  assign psq131 = sbd ? xs[131] : qs131;
  assign psq132 = sbd ? xs[132] : qs132;
  assign psq133 = sbd ? xs[133] : qs133;
  assign psq134 = sbd ? xs[134] : qs134;
  assign psq135 = sbd ? xs[135] : qs135;
  assign psq136 = sbd ? xs[136] : qs136;
  assign psq137 = sbd ? xs[137] : qs137;
  assign psq138 = sbd ? xs[138] : qs138;
  assign psq139 = sbd ? xs[139] : qs139;
  assign psq140 = sbd ? xs[140] : qs140;
  assign psq141 = sbd ? xs[141] : qs141;
  assign psq142 = sbd ? xs[142] : qs142;
  assign psq143 = sbd ? xs[143] : qs143;
  assign psq144 = sbd ? xs[144] : qs144;
  assign psq145 = sbd ? xs[145] : qs145;
  assign psq146 = sbd ? xs[146] : qs146;
  assign psq147 = sbd ? xs[147] : qs147;
  assign psq148 = sbd ? xs[148] : qs148;
  assign psq149 = sbd ? xs[149] : qs149;
  assign psq150 = sbd ? xs[150] : qs150;
  assign psq151 = sbd ? xs[151] : qs151;
  assign psq152 = sbd ? xs[152] : qs152;
  assign psq153 = sbd ? xs[153] : qs153;
  assign psq154 = sbd ? xs[154] : qs154;
  assign psq155 = sbd ? xs[155] : qs155;
  assign psq156 = sbd ? xs[156] : qs156;
  assign psq157 = sbd ? xs[157] : qs157;
  assign psq158 = sbd ? xs[158] : qs158;
  assign psq159 = sbd ? xs[159] : qs159;
  assign psq160 = sbd ? xs[160] : qs160;
  assign psq161 = sbd ? xs[161] : qs161;
  assign psq162 = sbd ? xs[162] : qs162;
  assign psq163 = sbd ? xs[163] : qs163;
  assign psq164 = sbd ? xs[164] : qs164;
  assign psq165 = sbd ? xs[165] : qs165;
  assign psq166 = sbd ? xs[166] : qs166;
  assign psq167 = sbd ? xs[167] : qs167;
  assign psq168 = sbd ? xs[168] : qs168;
  assign psq169 = sbd ? xs[169] : qs169;
  assign psq170 = sbd ? xs[170] : qs170;
  assign psq171 = sbd ? xs[171] : qs171;
  assign psq172 = sbd ? xs[172] : qs172;
  assign psq173 = sbd ? xs[173] : qs173;
  assign psq174 = sbd ? xs[174] : qs174;
  assign psq175 = sbd ? xs[175] : qs175;
  assign psq176 = sbd ? xs[176] : qs176;
  assign psq177 = sbd ? xs[177] : qs177;
  assign psq178 = sbd ? xs[178] : qs178;
  assign psq179 = sbd ? xs[179] : qs179;
  assign psq180 = sbd ? xs[180] : qs180;
  assign psq181 = sbd ? xs[181] : qs181;
  assign psq182 = sbd ? xs[182] : qs182;
  assign psq183 = sbd ? xs[183] : qs183;
  assign psr0 = sad ? psq0 : ys0_o;
  assign psr1 = sad ? psq1 : ys1_o;
  assign psr2 = sad ? psq2 : ys2_o;
  assign psr3 = sad ? psq3 : ys3_o;
  assign psr4 = sad ? psq4 : ys4_o;
  assign psr5 = sad ? psq5 : ys5_o;
  assign psr6 = sad ? psq6 : ys6_o;
  assign psr7 = sad ? psq7 : ys7_o;
  assign psr8 = sad ? psq8 : ys8_o;
  assign psr9 = sad ? psq9 : ys9_o;
  assign psr10 = sad ? psq10 : ys10_o;
  assign psr11 = sad ? psq11 : ys11_o;
  assign psr12 = sad ? psq12 : ys12_o;
  assign psr13 = sad ? psq13 : ys13_o;
  assign psr14 = sad ? psq14 : ys14_o;
  assign psr15 = sad ? psq15 : ys15_o;
  assign psr16 = sad ? psq16 : ys16_o;
  assign psr17 = sad ? psq17 : ys17_o;
  assign psr18 = sad ? psq18 : ys18_o;
  assign psr19 = sad ? psq19 : ys19_o;
  assign psr20 = sad ? psq20 : ys20_o;
  assign psr21 = sad ? psq21 : ys21_o;
  assign psr22 = sad ? psq22 : ys22_o;
  assign psr23 = sad ? psq23 : ys23_o;
  assign psr24 = sad ? psq24 : ys24_o;
  assign psr25 = sad ? psq25 : ys25_o;
  assign psr26 = sad ? psq26 : ys26_o;
  assign psr27 = sad ? psq27 : ys27_o;
  assign psr28 = sad ? psq28 : ys28_o;
  assign psr29 = sad ? psq29 : ys29_o;
  assign psr30 = sad ? psq30 : ys30_o;
  assign psr31 = sad ? psq31 : ys31_o;
  assign psr32 = sad ? psq32 : ys32_o;
  assign psr33 = sad ? psq33 : ys33_o;
  assign psr34 = sad ? psq34 : ys34_o;
  assign psr35 = sad ? psq35 : ys35_o;
  assign psr36 = sad ? psq36 : ys36_o;
  assign psr37 = sad ? psq37 : ys37_o;
  assign psr38 = sad ? psq38 : ys38_o;
  assign psr39 = sad ? psq39 : ys39_o;
  assign psr40 = sad ? psq40 : ys40_o;
  assign psr41 = sad ? psq41 : ys41_o;
  assign psr42 = sad ? psq42 : ys42_o;
  assign psr43 = sad ? psq43 : ys43_o;
  assign psr44 = sad ? psq44 : ys44_o;
  assign psr45 = sad ? psq45 : ys45_o;
  assign psr46 = sad ? psq46 : ys46_o;
  assign psr47 = sad ? psq47 : ys47_o;
  assign psr48 = sad ? psq48 : ys48_o;
  assign psr49 = sad ? psq49 : ys49_o;
  assign psr50 = sad ? psq50 : ys50_o;
  assign psr51 = sad ? psq51 : ys51_o;
  assign psr52 = sad ? psq52 : ys52_o;
  assign psr53 = sad ? psq53 : ys53_o;
  assign psr54 = sad ? psq54 : ys54_o;
  assign psr55 = sad ? psq55 : ys55_o;
  assign psr56 = sad ? psq56 : ys56_o;
  assign psr57 = sad ? psq57 : ys57_o;
  assign psr58 = sad ? psq58 : ys58_o;
  assign psr59 = sad ? psq59 : ys59_o;
  assign psr60 = sad ? psq60 : ys60_o;
  assign psr61 = sad ? psq61 : ys61_o;
  assign psr62 = sad ? psq62 : ys62_o;
  assign psr63 = sad ? psq63 : ys63_o;
  assign psr64 = sad ? psq64 : ys64_o;
  assign psr65 = sad ? psq65 : ys65_o;
  assign psr66 = sad ? psq66 : ys66_o;
  assign psr67 = sad ? psq67 : ys67_o;
  assign psr68 = sad ? psq68 : ys68_o;
  assign psr69 = sad ? psq69 : ys69_o;
  assign psr70 = sad ? psq70 : ys70_o;
  assign psr71 = sad ? psq71 : ys71_o;
  assign psr72 = sad ? psq72 : ys72_o;
  assign psr73 = sad ? psq73 : ys73_o;
  assign psr74 = sad ? psq74 : ys74_o;
  assign psr75 = sad ? psq75 : ys75_o;
  assign psr76 = sad ? psq76 : ys76_o;
  assign psr77 = sad ? psq77 : ys77_o;
  assign psr78 = sad ? psq78 : ys78_o;
  assign psr79 = sad ? psq79 : ys79_o;
  assign psr80 = sad ? psq80 : ys80_o;
  assign psr81 = sad ? psq81 : ys81_o;
  assign psr82 = sad ? psq82 : ys82_o;
  assign psr83 = sad ? psq83 : ys83_o;
  assign psr84 = sad ? psq84 : ys84_o;
  assign psr85 = sad ? psq85 : ys85_o;
  assign psr86 = sad ? psq86 : ys86_o;
  assign psr87 = sad ? psq87 : ys87_o;
  assign psr88 = sad ? psq88 : ys88_o;
  assign psr89 = sad ? psq89 : ys89_o;
  assign psr90 = sad ? psq90 : ys90_o;
  assign psr91 = sad ? psq91 : ys91_o;
  assign psr92 = sad ? psq92 : ys92_o;
  assign psr93 = sad ? psq93 : ys93_o;
  assign psr94 = sad ? psq94 : ys94_o;
  assign psr95 = sad ? psq95 : ys95_o;
  assign psr96 = sad ? psq96 : ys96_o;
  assign psr97 = sad ? psq97 : ys97_o;
  assign psr98 = sad ? psq98 : ys98_o;
  assign psr99 = sad ? psq99 : ys99_o;
  assign psr100 = sad ? psq100 : ys100_o;
  assign psr101 = sad ? psq101 : ys101_o;
  assign psr102 = sad ? psq102 : ys102_o;
  assign psr103 = sad ? psq103 : ys103_o;
  assign psr104 = sad ? psq104 : ys104_o;
  assign psr105 = sad ? psq105 : ys105_o;
  assign psr106 = sad ? psq106 : ys106_o;
  assign psr107 = sad ? psq107 : ys107_o;
  assign psr108 = sad ? psq108 : ys108_o;
  assign psr109 = sad ? psq109 : ys109_o;
  assign psr110 = sad ? psq110 : ys110_o;
  assign psr111 = sad ? psq111 : ys111_o;
  assign psr112 = sad ? psq112 : ys112_o;
  assign psr113 = sad ? psq113 : ys113_o;
  assign psr114 = sad ? psq114 : ys114_o;
  assign psr115 = sad ? psq115 : ys115_o;
  assign psr116 = sad ? psq116 : ys116_o;
  assign psr117 = sad ? psq117 : ys117_o;
  assign psr118 = sad ? psq118 : ys118_o;
  assign psr119 = sad ? psq119 : ys119_o;
  assign psr120 = sad ? psq120 : ys120_o;
  assign psr121 = sad ? psq121 : ys121_o;
  assign psr122 = sad ? psq122 : ys122_o;
  assign psr123 = sad ? psq123 : ys123_o;
  assign psr124 = sad ? psq124 : ys124_o;
  assign psr125 = sad ? psq125 : ys125_o;
  assign psr126 = sad ? psq126 : ys126_o;
  assign psr127 = sad ? psq127 : ys127_o;
  assign psr128 = sad ? psq128 : ys128_o;
  assign psr129 = sad ? psq129 : ys129_o;
  assign psr130 = sad ? psq130 : ys130_o;
  assign psr131 = sad ? psq131 : ys131_o;
  assign psr132 = sad ? psq132 : ys132_o;
  assign psr133 = sad ? psq133 : ys133_o;
  assign psr134 = sad ? psq134 : ys134_o;
  assign psr135 = sad ? psq135 : ys135_o;
  assign psr136 = sad ? psq136 : ys136_o;
  assign psr137 = sad ? psq137 : ys137_o;
  assign psr138 = sad ? psq138 : ys138_o;
  assign psr139 = sad ? psq139 : ys139_o;
  assign psr140 = sad ? psq140 : ys140_o;
  assign psr141 = sad ? psq141 : ys141_o;
  assign psr142 = sad ? psq142 : ys142_o;
  assign psr143 = sad ? psq143 : ys143_o;
  assign psr144 = sad ? psq144 : ys144_o;
  assign psr145 = sad ? psq145 : ys145_o;
  assign psr146 = sad ? psq146 : ys146_o;
  assign psr147 = sad ? psq147 : ys147_o;
  assign psr148 = sad ? psq148 : ys148_o;
  assign psr149 = sad ? psq149 : ys149_o;
  assign psr150 = sad ? psq150 : ys150_o;
  assign psr151 = sad ? psq151 : ys151_o;
  assign psr152 = sad ? psq152 : ys152_o;
  assign psr153 = sad ? psq153 : ys153_o;
  assign psr154 = sad ? psq154 : ys154_o;
  assign psr155 = sad ? psq155 : ys155_o;
  assign psr156 = sad ? psq156 : ys156_o;
  assign psr157 = sad ? psq157 : ys157_o;
  assign psr158 = sad ? psq158 : ys158_o;
  assign psr159 = sad ? psq159 : ys159_o;
  assign psr160 = sad ? psq160 : ys160_o;
  assign psr161 = sad ? psq161 : ys161_o;
  assign psr162 = sad ? psq162 : ys162_o;
  assign psr163 = sad ? psq163 : ys163_o;
  assign psr164 = sad ? psq164 : ys164_o;
  assign psr165 = sad ? psq165 : ys165_o;
  assign psr166 = sad ? psq166 : ys166_o;
  assign psr167 = sad ? psq167 : ys167_o;
  assign psr168 = sad ? psq168 : ys168_o;
  assign psr169 = sad ? psq169 : ys169_o;
  assign psr170 = sad ? psq170 : ys170_o;
  assign psr171 = sad ? psq171 : ys171_o;
  assign psr172 = sad ? psq172 : ys172_o;
  assign psr173 = sad ? psq173 : ys173_o;
  assign psr174 = sad ? psq174 : ys174_o;
  assign psr175 = sad ? psq175 : ys175_o;
  assign psr176 = sad ? psq176 : ys176_o;
  assign psr177 = sad ? psq177 : ys177_o;
  assign psr178 = sad ? psq178 : ys178_o;
  assign psr179 = sad ? psq179 : ys179_o;
  assign psr180 = sad ? psq180 : ys180_o;
  assign psr181 = sad ? psq181 : ys181_o;
  assign psr182 = sad ? psq182 : ys182_o;
  assign psr183 = sad ? psq183 : ys183_o;
  assign qc0 = multm_qsp0 & multm_compress_nsd;
  assign qc1 = multm_compress_add3b_maj3b_or3b_wx0 | multm_compress_add3b_maj3b_xy0;
  assign qc2 = multm_qsp2 & multm_qcp1;
  assign qc3 = multm_compress_add3b_maj3b_or3b_wx2 | multm_compress_add3b_maj3b_xy2;
  assign qc4 = multm_compress_add3b_maj3b_or3b_wx3 | multm_compress_add3b_maj3b_xy3;
  assign qc5 = multm_compress_add3b_maj3b_or3b_wx4 | multm_compress_add3b_maj3b_xy4;
  assign qc6 = multm_compress_add3b_maj3b_or3b_wx5 | multm_compress_add3b_maj3b_xy5;
  assign qc7 = multm_qsp7 & multm_qcp6;
  assign qc8 = multm_qsp8 & multm_qcp7;
  assign qc9 = multm_compress_add3b_maj3b_or3b_wx8 | multm_compress_add3b_maj3b_xy8;
  assign qc10 = multm_compress_add3b_maj3b_or3b_wx9 | multm_compress_add3b_maj3b_xy9;
  assign qc11 = multm_compress_add3b_maj3b_or3b_wx10 | multm_compress_add3b_maj3b_xy10;
  assign qc12 = multm_compress_add3b_maj3b_or3b_wx11 | multm_compress_add3b_maj3b_xy11;
  assign qc13 = multm_compress_add3b_maj3b_or3b_wx12 | multm_compress_add3b_maj3b_xy12;
  assign qc14 = multm_compress_add3b_maj3b_or3b_wx13 | multm_compress_add3b_maj3b_xy13;
  assign qc15 = multm_compress_add3b_maj3b_or3b_wx14 | multm_compress_add3b_maj3b_xy14;
  assign qc16 = multm_compress_add3b_maj3b_or3b_wx15 | multm_compress_add3b_maj3b_xy15;
  assign qc17 = multm_compress_add3b_maj3b_or3b_wx16 | multm_compress_add3b_maj3b_xy16;
  assign qc18 = multm_compress_add3b_maj3b_or3b_wx17 | multm_compress_add3b_maj3b_xy17;
  assign qc19 = multm_compress_add3b_maj3b_or3b_wx18 | multm_compress_add3b_maj3b_xy18;
  assign qc20 = multm_compress_add3b_maj3b_or3b_wx19 | multm_compress_add3b_maj3b_xy19;
  assign qc21 = multm_compress_add3b_maj3b_or3b_wx20 | multm_compress_add3b_maj3b_xy20;
  assign qc22 = multm_compress_add3b_maj3b_or3b_wx21 | multm_compress_add3b_maj3b_xy21;
  assign qc23 = multm_compress_add3b_maj3b_or3b_wx22 | multm_compress_add3b_maj3b_xy22;
  assign qc24 = multm_compress_add3b_maj3b_or3b_wx23 | multm_compress_add3b_maj3b_xy23;
  assign qc25 = multm_qsp25 & multm_qcp24;
  assign qc26 = multm_compress_add3b_maj3b_or3b_wx25 | multm_compress_add3b_maj3b_xy25;
  assign qc27 = multm_compress_add3b_maj3b_or3b_wx26 | multm_compress_add3b_maj3b_xy26;
  assign qc28 = multm_compress_add3b_maj3b_or3b_wx27 | multm_compress_add3b_maj3b_xy27;
  assign qc29 = multm_compress_add3b_maj3b_or3b_wx28 | multm_compress_add3b_maj3b_xy28;
  assign qc30 = multm_compress_add3b_maj3b_or3b_wx29 | multm_compress_add3b_maj3b_xy29;
  assign qc31 = multm_compress_add3b_maj3b_or3b_wx30 | multm_compress_add3b_maj3b_xy30;
  assign qc32 = multm_compress_add3b_maj3b_or3b_wx31 | multm_compress_add3b_maj3b_xy31;
  assign qc33 = multm_compress_add3b_maj3b_or3b_wx32 | multm_compress_add3b_maj3b_xy32;
  assign qc34 = multm_compress_add3b_maj3b_or3b_wx33 | multm_compress_add3b_maj3b_xy33;
  assign qc35 = multm_compress_add3b_maj3b_or3b_wx34 | multm_compress_add3b_maj3b_xy34;
  assign qc36 = multm_compress_add3b_maj3b_or3b_wx35 | multm_compress_add3b_maj3b_xy35;
  assign qc37 = multm_compress_add3b_maj3b_or3b_wx36 | multm_compress_add3b_maj3b_xy36;
  assign qc38 = multm_compress_add3b_maj3b_or3b_wx37 | multm_compress_add3b_maj3b_xy37;
  assign qc39 = multm_compress_add3b_maj3b_or3b_wx38 | multm_compress_add3b_maj3b_xy38;
  assign qc40 = multm_compress_add3b_maj3b_or3b_wx39 | multm_compress_add3b_maj3b_xy39;
  assign qc41 = multm_compress_add3b_maj3b_or3b_wx40 | multm_compress_add3b_maj3b_xy40;
  assign qc42 = multm_compress_add3b_maj3b_or3b_wx41 | multm_compress_add3b_maj3b_xy41;
  assign qc43 = multm_qsp43 & multm_qcp42;
  assign qc44 = multm_qsp44 & multm_qcp43;
  assign qc45 = multm_compress_add3b_maj3b_or3b_wx44 | multm_compress_add3b_maj3b_xy44;
  assign qc46 = multm_compress_add3b_maj3b_or3b_wx45 | multm_compress_add3b_maj3b_xy45;
  assign qc47 = multm_compress_add3b_maj3b_or3b_wx46 | multm_compress_add3b_maj3b_xy46;
  assign qc48 = multm_compress_add3b_maj3b_or3b_wx47 | multm_compress_add3b_maj3b_xy47;
  assign qc49 = multm_compress_add3b_maj3b_or3b_wx48 | multm_compress_add3b_maj3b_xy48;
  assign qc50 = multm_compress_add3b_maj3b_or3b_wx49 | multm_compress_add3b_maj3b_xy49;
  assign qc51 = multm_compress_add3b_maj3b_or3b_wx50 | multm_compress_add3b_maj3b_xy50;
  assign qc52 = multm_compress_add3b_maj3b_or3b_wx51 | multm_compress_add3b_maj3b_xy51;
  assign qc53 = multm_compress_add3b_maj3b_or3b_wx52 | multm_compress_add3b_maj3b_xy52;
  assign qc54 = multm_qsp54 & multm_qcp53;
  assign qc55 = multm_qsp55 & multm_qcp54;
  assign qc56 = multm_qsp56 & multm_qcp55;
  assign qc57 = multm_compress_add3b_maj3b_or3b_wx56 | multm_compress_add3b_maj3b_xy56;
  assign qc58 = multm_compress_add3b_maj3b_or3b_wx57 | multm_compress_add3b_maj3b_xy57;
  assign qc59 = multm_compress_add3b_maj3b_or3b_wx58 | multm_compress_add3b_maj3b_xy58;
  assign qc60 = multm_compress_add3b_maj3b_or3b_wx59 | multm_compress_add3b_maj3b_xy59;
  assign qc61 = multm_compress_add3b_maj3b_or3b_wx60 | multm_compress_add3b_maj3b_xy60;
  assign qc62 = multm_compress_add3b_maj3b_or3b_wx61 | multm_compress_add3b_maj3b_xy61;
  assign qc63 = multm_compress_add3b_maj3b_or3b_wx62 | multm_compress_add3b_maj3b_xy62;
  assign qc64 = multm_compress_add3b_maj3b_or3b_wx63 | multm_compress_add3b_maj3b_xy63;
  assign qc65 = multm_compress_add3b_maj3b_or3b_wx64 | multm_compress_add3b_maj3b_xy64;
  assign qc66 = multm_compress_add3b_maj3b_or3b_wx65 | multm_compress_add3b_maj3b_xy65;
  assign qc67 = multm_compress_add3b_maj3b_or3b_wx66 | multm_compress_add3b_maj3b_xy66;
  assign qc68 = multm_compress_add3b_maj3b_or3b_wx67 | multm_compress_add3b_maj3b_xy67;
  assign qc69 = multm_compress_add3b_maj3b_or3b_wx68 | multm_compress_add3b_maj3b_xy68;
  assign qc70 = multm_compress_add3b_maj3b_or3b_wx69 | multm_compress_add3b_maj3b_xy69;
  assign qc71 = multm_compress_add3b_maj3b_or3b_wx70 | multm_compress_add3b_maj3b_xy70;
  assign qc72 = multm_compress_add3b_maj3b_or3b_wx71 | multm_compress_add3b_maj3b_xy71;
  assign qc73 = multm_compress_add3b_maj3b_or3b_wx72 | multm_compress_add3b_maj3b_xy72;
  assign qc74 = multm_compress_add3b_maj3b_or3b_wx73 | multm_compress_add3b_maj3b_xy73;
  assign qc75 = multm_qsp75 & multm_qcp74;
  assign qc76 = multm_compress_add3b_maj3b_or3b_wx75 | multm_compress_add3b_maj3b_xy75;
  assign qc77 = multm_compress_add3b_maj3b_or3b_wx76 | multm_compress_add3b_maj3b_xy76;
  assign qc78 = multm_compress_add3b_maj3b_or3b_wx77 | multm_compress_add3b_maj3b_xy77;
  assign qc79 = multm_compress_add3b_maj3b_or3b_wx78 | multm_compress_add3b_maj3b_xy78;
  assign qc80 = multm_compress_add3b_maj3b_or3b_wx79 | multm_compress_add3b_maj3b_xy79;
  assign qc81 = multm_compress_add3b_maj3b_or3b_wx80 | multm_compress_add3b_maj3b_xy80;
  assign qc82 = multm_compress_add3b_maj3b_or3b_wx81 | multm_compress_add3b_maj3b_xy81;
  assign qc83 = multm_compress_add3b_maj3b_or3b_wx82 | multm_compress_add3b_maj3b_xy82;
  assign qc84 = multm_compress_add3b_maj3b_or3b_wx83 | multm_compress_add3b_maj3b_xy83;
  assign qc85 = multm_compress_add3b_maj3b_or3b_wx84 | multm_compress_add3b_maj3b_xy84;
  assign qc86 = multm_compress_add3b_maj3b_or3b_wx85 | multm_compress_add3b_maj3b_xy85;
  assign qc87 = multm_compress_add3b_maj3b_or3b_wx86 | multm_compress_add3b_maj3b_xy86;
  assign qc88 = multm_compress_add3b_maj3b_or3b_wx87 | multm_compress_add3b_maj3b_xy87;
  assign qc89 = multm_compress_add3b_maj3b_or3b_wx88 | multm_compress_add3b_maj3b_xy88;
  assign qc90 = multm_compress_add3b_maj3b_or3b_wx89 | multm_compress_add3b_maj3b_xy89;
  assign qc91 = multm_compress_add3b_maj3b_or3b_wx90 | multm_compress_add3b_maj3b_xy90;
  assign qc92 = multm_compress_add3b_maj3b_or3b_wx91 | multm_compress_add3b_maj3b_xy91;
  assign qc93 = multm_compress_add3b_maj3b_or3b_wx92 | multm_compress_add3b_maj3b_xy92;
  assign qc94 = multm_compress_add3b_maj3b_or3b_wx93 | multm_compress_add3b_maj3b_xy93;
  assign qc95 = multm_compress_add3b_maj3b_or3b_wx94 | multm_compress_add3b_maj3b_xy94;
  assign qc96 = multm_compress_add3b_maj3b_or3b_wx95 | multm_compress_add3b_maj3b_xy95;
  assign qc97 = multm_compress_add3b_maj3b_or3b_wx96 | multm_compress_add3b_maj3b_xy96;
  assign qc98 = multm_compress_add3b_maj3b_or3b_wx97 | multm_compress_add3b_maj3b_xy97;
  assign qc99 = multm_compress_add3b_maj3b_or3b_wx98 | multm_compress_add3b_maj3b_xy98;
  assign qc100 = multm_compress_add3b_maj3b_or3b_wx99 | multm_compress_add3b_maj3b_xy99;
  assign qc101 = multm_compress_add3b_maj3b_or3b_wx100 | multm_compress_add3b_maj3b_xy100;
  assign qc102 = multm_qsp102 & multm_qcp101;
  assign qc103 = multm_qsp103 & multm_qcp102;
  assign qc104 = multm_compress_add3b_maj3b_or3b_wx103 | multm_compress_add3b_maj3b_xy103;
  assign qc105 = multm_compress_add3b_maj3b_or3b_wx104 | multm_compress_add3b_maj3b_xy104;
  assign qc106 = multm_qsp106 & multm_qcp105;
  assign qc107 = multm_compress_add3b_maj3b_or3b_wx106 | multm_compress_add3b_maj3b_xy106;
  assign qc108 = multm_compress_add3b_maj3b_or3b_wx107 | multm_compress_add3b_maj3b_xy107;
  assign qc109 = multm_qsp109 & multm_qcp108;
  assign qc110 = multm_qsp110 & multm_qcp109;
  assign qc111 = multm_qsp111 & multm_qcp110;
  assign qc112 = multm_compress_add3b_maj3b_or3b_wx111 | multm_compress_add3b_maj3b_xy111;
  assign qc113 = multm_compress_add3b_maj3b_or3b_wx112 | multm_compress_add3b_maj3b_xy112;
  assign qc114 = multm_compress_add3b_maj3b_or3b_wx113 | multm_compress_add3b_maj3b_xy113;
  assign qc115 = multm_compress_add3b_maj3b_or3b_wx114 | multm_compress_add3b_maj3b_xy114;
  assign qc116 = multm_compress_add3b_maj3b_or3b_wx115 | multm_compress_add3b_maj3b_xy115;
  assign qc117 = multm_compress_add3b_maj3b_or3b_wx116 | multm_compress_add3b_maj3b_xy116;
  assign qc118 = multm_compress_add3b_maj3b_or3b_wx117 | multm_compress_add3b_maj3b_xy117;
  assign qc119 = multm_compress_add3b_maj3b_or3b_wx118 | multm_compress_add3b_maj3b_xy118;
  assign qc120 = multm_qsp120 & multm_qcp119;
  assign qc121 = multm_qsp121 & multm_qcp120;
  assign qc122 = multm_qsp122 & multm_qcp121;
  assign qc123 = multm_qsp123 & multm_qcp122;
  assign qc124 = multm_qsp124 & multm_qcp123;
  assign qc125 = multm_compress_add3b_maj3b_or3b_wx124 | multm_compress_add3b_maj3b_xy124;
  assign qc126 = multm_compress_add3b_maj3b_or3b_wx125 | multm_compress_add3b_maj3b_xy125;
  assign qc127 = multm_compress_add3b_maj3b_or3b_wx126 | multm_compress_add3b_maj3b_xy126;
  assign qc128 = multm_compress_add3b_maj3b_or3b_wx127 | multm_compress_add3b_maj3b_xy127;
  assign qc129 = multm_compress_add3b_maj3b_or3b_wx128 | multm_compress_add3b_maj3b_xy128;
  assign qc130 = multm_compress_add3b_maj3b_or3b_wx129 | multm_compress_add3b_maj3b_xy129;
  assign qc131 = multm_compress_add3b_maj3b_or3b_wx130 | multm_compress_add3b_maj3b_xy130;
  assign qc132 = multm_compress_add3b_maj3b_or3b_wx131 | multm_compress_add3b_maj3b_xy131;
  assign qc133 = multm_compress_add3b_maj3b_or3b_wx132 | multm_compress_add3b_maj3b_xy132;
  assign qc134 = multm_compress_add3b_maj3b_or3b_wx133 | multm_compress_add3b_maj3b_xy133;
  assign qc135 = multm_compress_add3b_maj3b_or3b_wx134 | multm_compress_add3b_maj3b_xy134;
  assign qc136 = multm_compress_add3b_maj3b_or3b_wx135 | multm_compress_add3b_maj3b_xy135;
  assign qc137 = multm_compress_add3b_maj3b_or3b_wx136 | multm_compress_add3b_maj3b_xy136;
  assign qc138 = multm_compress_add3b_maj3b_or3b_wx137 | multm_compress_add3b_maj3b_xy137;
  assign qc139 = multm_compress_add3b_maj3b_or3b_wx138 | multm_compress_add3b_maj3b_xy138;
  assign qc140 = multm_compress_add3b_maj3b_or3b_wx139 | multm_compress_add3b_maj3b_xy139;
  assign qc141 = multm_compress_add3b_maj3b_or3b_wx140 | multm_compress_add3b_maj3b_xy140;
  assign qc142 = multm_compress_add3b_maj3b_or3b_wx141 | multm_compress_add3b_maj3b_xy141;
  assign qc143 = multm_qsp143 & multm_qcp142;
  assign qc144 = multm_qsp144 & multm_qcp143;
  assign qc145 = multm_qsp145 & multm_qcp144;
  assign qc146 = multm_compress_add3b_maj3b_or3b_wx145 | multm_compress_add3b_maj3b_xy145;
  assign qc147 = multm_compress_add3b_maj3b_or3b_wx146 | multm_compress_add3b_maj3b_xy146;
  assign qc148 = multm_compress_add3b_maj3b_or3b_wx147 | multm_compress_add3b_maj3b_xy147;
  assign qc149 = multm_compress_add3b_maj3b_or3b_wx148 | multm_compress_add3b_maj3b_xy148;
  assign qc150 = multm_compress_add3b_maj3b_or3b_wx149 | multm_compress_add3b_maj3b_xy149;
  assign qc151 = multm_compress_add3b_maj3b_or3b_wx150 | multm_compress_add3b_maj3b_xy150;
  assign qc152 = multm_compress_add3b_maj3b_or3b_wx151 | multm_compress_add3b_maj3b_xy151;
  assign qc153 = multm_qsp153 & multm_qcp152;
  assign qc154 = multm_qsp154 & multm_qcp153;
  assign qc155 = multm_compress_add3b_maj3b_or3b_wx154 | multm_compress_add3b_maj3b_xy154;
  assign qc156 = multm_compress_add3b_maj3b_or3b_wx155 | multm_compress_add3b_maj3b_xy155;
  assign qc157 = multm_qsp157 & multm_qcp156;
  assign qc158 = multm_qsp158 & multm_qcp157;
  assign qc159 = multm_qsp159 & multm_qcp158;
  assign qc160 = multm_qsp160 & multm_qcp159;
  assign qc161 = multm_qsp161 & multm_qcp160;
  assign qc162 = multm_compress_add3b_maj3b_or3b_wx161 | multm_compress_add3b_maj3b_xy161;
  assign qc163 = multm_compress_add3b_maj3b_or3b_wx162 | multm_compress_add3b_maj3b_xy162;
  assign qc164 = multm_compress_add3b_maj3b_or3b_wx163 | multm_compress_add3b_maj3b_xy163;
  assign qc165 = multm_compress_add3b_maj3b_or3b_wx164 | multm_compress_add3b_maj3b_xy164;
  assign qc166 = multm_compress_add3b_maj3b_or3b_wx165 | multm_compress_add3b_maj3b_xy165;
  assign qc167 = multm_compress_add3b_maj3b_or3b_wx166 | multm_compress_add3b_maj3b_xy166;
  assign qc168 = multm_compress_add3b_maj3b_or3b_wx167 | multm_compress_add3b_maj3b_xy167;
  assign qc169 = multm_compress_add3b_maj3b_or3b_wx168 | multm_compress_add3b_maj3b_xy168;
  assign qc170 = multm_compress_add3b_maj3b_or3b_wx169 | multm_compress_add3b_maj3b_xy169;
  assign qc171 = multm_compress_add3b_maj3b_or3b_wx170 | multm_compress_add3b_maj3b_xy170;
  assign qc172 = multm_compress_add3b_maj3b_or3b_wx171 | multm_compress_add3b_maj3b_xy171;
  assign qc173 = multm_compress_add3b_maj3b_or3b_wx172 | multm_compress_add3b_maj3b_xy172;
  assign qc174 = multm_qsp174 & multm_qcp173;
  assign qc175 = multm_qsp175 & multm_qcp174;
  assign qc176 = multm_qsp176 & multm_qcp175;
  assign qc177 = multm_compress_add3b_maj3b_or3b_wx176 | multm_compress_add3b_maj3b_xy176;
  assign qc178 = multm_compress_add3b_maj3b_or3b_wx177 | multm_compress_add3b_maj3b_xy177;
  assign qc179 = multm_compress_add3b_maj3b_or3b_wx178 | multm_compress_add3b_maj3b_xy178;
  assign qc180 = multm_compress_add3b_maj3b_or3b_wx179 | multm_compress_add3b_maj3b_xy179;
  assign qc181 = multm_compress_add3b_maj3b_or3b_wx180 | multm_compress_add3b_maj3b_xy180;
  assign qc182 = multm_compress_add3b_maj3b_or3b_wx181 | multm_compress_add3b_maj3b_xy181;
  assign qc183 = multm_compress_add3b_maj3b_or3b_wx182 | multm_compress_add3b_maj3b_xy182;
  assign qs0 = multm_qsp0 ^ multm_compress_nsd;
  assign qs1 = multm_compress_add3b_xor3b_wx0 ^ multm_compress_ncd;
  assign qs2 = multm_qsp2 ^ multm_qcp1;
  assign qs3 = multm_compress_add3b_xor3b_wx2 ^ multm_compress_nsd;
  assign qs4 = multm_compress_add3b_xor3b_wx3 ^ multm_compress_rn4;
  assign qs5 = multm_compress_add3b_xor3b_wx4 ^ multm_compress_rn5;
  assign qs6 = multm_compress_add3b_xor3b_wx5 ^ multm_compress_rn6;
  assign qs7 = multm_qsp7 ^ multm_qcp6;
  assign qs8 = multm_qsp8 ^ multm_qcp7;
  assign qs9 = multm_compress_add3b_xor3b_wx8 ^ multm_compress_nsd;
  assign qs10 = multm_compress_add3b_xor3b_wx9 ^ multm_compress_rn4;
  assign qs11 = multm_compress_add3b_xor3b_wx10 ^ multm_compress_rn5;
  assign qs12 = multm_compress_add3b_xor3b_wx11 ^ multm_compress_rn20;
  assign qs13 = multm_compress_add3b_xor3b_wx12 ^ multm_compress_rn5;
  assign qs14 = multm_compress_add3b_xor3b_wx13 ^ multm_compress_rn20;
  assign qs15 = multm_compress_add3b_xor3b_wx14 ^ multm_compress_rn15;
  assign qs16 = multm_compress_add3b_xor3b_wx15 ^ multm_compress_rn15;
  assign qs17 = multm_compress_add3b_xor3b_wx16 ^ multm_compress_rn15;
  assign qs18 = multm_compress_add3b_xor3b_wx17 ^ multm_compress_rn15;
  assign qs19 = multm_compress_add3b_xor3b_wx18 ^ multm_compress_rn5;
  assign qs20 = multm_compress_add3b_xor3b_wx19 ^ multm_compress_rn20;
  assign qs21 = multm_compress_add3b_xor3b_wx20 ^ multm_compress_rn5;
  assign qs22 = multm_compress_add3b_xor3b_wx21 ^ multm_compress_rn20;
  assign qs23 = multm_compress_add3b_xor3b_wx22 ^ multm_compress_rn5;
  assign qs24 = multm_compress_add3b_xor3b_wx23 ^ multm_compress_rn6;
  assign qs25 = multm_qsp25 ^ multm_qcp24;
  assign qs26 = multm_compress_add3b_xor3b_wx25 ^ multm_compress_nsd;
  assign qs27 = multm_compress_add3b_xor3b_wx26 ^ multm_compress_rn4;
  assign qs28 = multm_compress_add3b_xor3b_wx27 ^ multm_compress_rn15;
  assign qs29 = multm_compress_add3b_xor3b_wx28 ^ multm_compress_rn5;
  assign qs30 = multm_compress_add3b_xor3b_wx29 ^ multm_compress_rn20;
  assign qs31 = multm_compress_add3b_xor3b_wx30 ^ multm_compress_rn5;
  assign qs32 = multm_compress_add3b_xor3b_wx31 ^ multm_compress_rn20;
  assign qs33 = multm_compress_add3b_xor3b_wx32 ^ multm_compress_rn5;
  assign qs34 = multm_compress_add3b_xor3b_wx33 ^ multm_compress_rn20;
  assign qs35 = multm_compress_add3b_xor3b_wx34 ^ multm_compress_rn5;
  assign qs36 = multm_compress_add3b_xor3b_wx35 ^ multm_compress_rn20;
  assign qs37 = multm_compress_add3b_xor3b_wx36 ^ multm_compress_rn15;
  assign qs38 = multm_compress_add3b_xor3b_wx37 ^ multm_compress_rn5;
  assign qs39 = multm_compress_add3b_xor3b_wx38 ^ multm_compress_rn20;
  assign qs40 = multm_compress_add3b_xor3b_wx39 ^ multm_compress_rn15;
  assign qs41 = multm_compress_add3b_xor3b_wx40 ^ multm_compress_rn5;
  assign qs42 = multm_compress_add3b_xor3b_wx41 ^ multm_compress_rn6;
  assign qs43 = multm_qsp43 ^ multm_qcp42;
  assign qs44 = multm_qsp44 ^ multm_qcp43;
  assign qs45 = multm_compress_add3b_xor3b_wx44 ^ multm_compress_nsd;
  assign qs46 = multm_compress_add3b_xor3b_wx45 ^ multm_compress_rn4;
  assign qs47 = multm_compress_add3b_xor3b_wx46 ^ multm_compress_rn15;
  assign qs48 = multm_compress_add3b_xor3b_wx47 ^ multm_compress_rn5;
  assign qs49 = multm_compress_add3b_xor3b_wx48 ^ multm_compress_rn6;
  assign qs50 = multm_compress_add3b_xor3b_wx49 ^ multm_compress_nsd;
  assign qs51 = multm_compress_add3b_xor3b_wx50 ^ multm_compress_rn4;
  assign qs52 = multm_compress_add3b_xor3b_wx51 ^ multm_compress_rn5;
  assign qs53 = multm_compress_add3b_xor3b_wx52 ^ multm_compress_rn6;
  assign qs54 = multm_qsp54 ^ multm_qcp53;
  assign qs55 = multm_qsp55 ^ multm_qcp54;
  assign qs56 = multm_qsp56 ^ multm_qcp55;
  assign qs57 = multm_compress_add3b_xor3b_wx56 ^ multm_compress_nsd;
  assign qs58 = multm_compress_add3b_xor3b_wx57 ^ multm_compress_ncd;
  assign qs59 = multm_compress_add3b_xor3b_wx58 ^ multm_compress_nsd;
  assign qs60 = multm_compress_add3b_xor3b_wx59 ^ multm_compress_rn4;
  assign qs61 = multm_compress_add3b_xor3b_wx60 ^ multm_compress_rn15;
  assign qs62 = multm_compress_add3b_xor3b_wx61 ^ multm_compress_rn15;
  assign qs63 = multm_compress_add3b_xor3b_wx62 ^ multm_compress_rn5;
  assign qs64 = multm_compress_add3b_xor3b_wx63 ^ multm_compress_rn20;
  assign qs65 = multm_compress_add3b_xor3b_wx64 ^ multm_compress_rn15;
  assign qs66 = multm_compress_add3b_xor3b_wx65 ^ multm_compress_rn15;
  assign qs67 = multm_compress_add3b_xor3b_wx66 ^ multm_compress_rn5;
  assign qs68 = multm_compress_add3b_xor3b_wx67 ^ multm_compress_rn20;
  assign qs69 = multm_compress_add3b_xor3b_wx68 ^ multm_compress_rn5;
  assign qs70 = multm_compress_add3b_xor3b_wx69 ^ multm_compress_rn6;
  assign qs71 = multm_compress_add3b_xor3b_wx70 ^ multm_compress_nsd;
  assign qs72 = multm_compress_add3b_xor3b_wx71 ^ multm_compress_ncd;
  assign qs73 = multm_compress_add3b_xor3b_wx72 ^ multm_compress_nsd;
  assign qs74 = multm_compress_add3b_xor3b_wx73 ^ multm_compress_ncd;
  assign qs75 = multm_qsp75 ^ multm_qcp74;
  assign qs76 = multm_compress_add3b_xor3b_wx75 ^ multm_compress_nsd;
  assign qs77 = multm_compress_add3b_xor3b_wx76 ^ multm_compress_rn4;
  assign qs78 = multm_compress_add3b_xor3b_wx77 ^ multm_compress_rn15;
  assign qs79 = multm_compress_add3b_xor3b_wx78 ^ multm_compress_rn15;
  assign qs80 = multm_compress_add3b_xor3b_wx79 ^ multm_compress_rn5;
  assign qs81 = multm_compress_add3b_xor3b_wx80 ^ multm_compress_rn6;
  assign qs82 = multm_compress_add3b_xor3b_wx81 ^ multm_compress_nsd;
  assign qs83 = multm_compress_add3b_xor3b_wx82 ^ multm_compress_ncd;
  assign qs84 = multm_compress_add3b_xor3b_wx83 ^ multm_compress_nsd;
  assign qs85 = multm_compress_add3b_xor3b_wx84 ^ multm_compress_rn4;
  assign qs86 = multm_compress_add3b_xor3b_wx85 ^ multm_compress_rn15;
  assign qs87 = multm_compress_add3b_xor3b_wx86 ^ multm_compress_rn5;
  assign qs88 = multm_compress_add3b_xor3b_wx87 ^ multm_compress_rn20;
  assign qs89 = multm_compress_add3b_xor3b_wx88 ^ multm_compress_rn5;
  assign qs90 = multm_compress_add3b_xor3b_wx89 ^ multm_compress_rn20;
  assign qs91 = multm_compress_add3b_xor3b_wx90 ^ multm_compress_rn5;
  assign qs92 = multm_compress_add3b_xor3b_wx91 ^ multm_compress_rn6;
  assign qs93 = multm_compress_add3b_xor3b_wx92 ^ multm_compress_nsd;
  assign qs94 = multm_compress_add3b_xor3b_wx93 ^ multm_compress_rn4;
  assign qs95 = multm_compress_add3b_xor3b_wx94 ^ multm_compress_rn15;
  assign qs96 = multm_compress_add3b_xor3b_wx95 ^ multm_compress_rn15;
  assign qs97 = multm_compress_add3b_xor3b_wx96 ^ multm_compress_rn5;
  assign qs98 = multm_compress_add3b_xor3b_wx97 ^ multm_compress_rn20;
  assign qs99 = multm_compress_add3b_xor3b_wx98 ^ multm_compress_rn15;
  assign qs100 = multm_compress_add3b_xor3b_wx99 ^ multm_compress_rn5;
  assign qs101 = multm_compress_add3b_xor3b_wx100 ^ multm_compress_rn6;
  assign qs102 = multm_qsp102 ^ multm_qcp101;
  assign qs103 = multm_qsp103 ^ multm_qcp102;
  assign qs104 = multm_compress_add3b_xor3b_wx103 ^ multm_compress_nsd;
  assign qs105 = multm_compress_add3b_xor3b_wx104 ^ multm_compress_ncd;
  assign qs106 = multm_qsp106 ^ multm_qcp105;
  assign qs107 = multm_compress_add3b_xor3b_wx106 ^ multm_compress_nsd;
  assign qs108 = multm_compress_add3b_xor3b_wx107 ^ multm_compress_ncd;
  assign qs109 = multm_qsp109 ^ multm_qcp108;
  assign qs110 = multm_qsp110 ^ multm_qcp109;
  assign qs111 = multm_qsp111 ^ multm_qcp110;
  assign qs112 = multm_compress_add3b_xor3b_wx111 ^ multm_compress_nsd;
  assign qs113 = multm_compress_add3b_xor3b_wx112 ^ multm_compress_ncd;
  assign qs114 = multm_compress_add3b_xor3b_wx113 ^ multm_compress_nsd;
  assign qs115 = multm_compress_add3b_xor3b_wx114 ^ multm_compress_ncd;
  assign qs116 = multm_compress_add3b_xor3b_wx115 ^ multm_compress_nsd;
  assign qs117 = multm_compress_add3b_xor3b_wx116 ^ multm_compress_rn4;
  assign qs118 = multm_compress_add3b_xor3b_wx117 ^ multm_compress_rn5;
  assign qs119 = multm_compress_add3b_xor3b_wx118 ^ multm_compress_rn6;
  assign qs120 = multm_qsp120 ^ multm_qcp119;
  assign qs121 = multm_qsp121 ^ multm_qcp120;
  assign qs122 = multm_qsp122 ^ multm_qcp121;
  assign qs123 = multm_qsp123 ^ multm_qcp122;
  assign qs124 = multm_qsp124 ^ multm_qcp123;
  assign qs125 = multm_compress_add3b_xor3b_wx124 ^ multm_compress_nsd;
  assign qs126 = multm_compress_add3b_xor3b_wx125 ^ multm_compress_rn4;
  assign qs127 = multm_compress_add3b_xor3b_wx126 ^ multm_compress_rn15;
  assign qs128 = multm_compress_add3b_xor3b_wx127 ^ multm_compress_rn15;
  assign qs129 = multm_compress_add3b_xor3b_wx128 ^ multm_compress_rn5;
  assign qs130 = multm_compress_add3b_xor3b_wx129 ^ multm_compress_rn20;
  assign qs131 = multm_compress_add3b_xor3b_wx130 ^ multm_compress_rn5;
  assign qs132 = multm_compress_add3b_xor3b_wx131 ^ multm_compress_rn20;
  assign qs133 = multm_compress_add3b_xor3b_wx132 ^ multm_compress_rn5;
  assign qs134 = multm_compress_add3b_xor3b_wx133 ^ multm_compress_rn20;
  assign qs135 = multm_compress_add3b_xor3b_wx134 ^ multm_compress_rn15;
  assign qs136 = multm_compress_add3b_xor3b_wx135 ^ multm_compress_rn5;
  assign qs137 = multm_compress_add3b_xor3b_wx136 ^ multm_compress_rn6;
  assign qs138 = multm_compress_add3b_xor3b_wx137 ^ multm_compress_nsd;
  assign qs139 = multm_compress_add3b_xor3b_wx138 ^ multm_compress_rn4;
  assign qs140 = multm_compress_add3b_xor3b_wx139 ^ multm_compress_rn15;
  assign qs141 = multm_compress_add3b_xor3b_wx140 ^ multm_compress_rn5;
  assign qs142 = multm_compress_add3b_xor3b_wx141 ^ multm_compress_rn6;
  assign qs143 = multm_qsp143 ^ multm_qcp142;
  assign qs144 = multm_qsp144 ^ multm_qcp143;
  assign qs145 = multm_qsp145 ^ multm_qcp144;
  assign qs146 = multm_compress_add3b_xor3b_wx145 ^ multm_compress_nsd;
  assign qs147 = multm_compress_add3b_xor3b_wx146 ^ multm_compress_rn4;
  assign qs148 = multm_compress_add3b_xor3b_wx147 ^ multm_compress_rn5;
  assign qs149 = multm_compress_add3b_xor3b_wx148 ^ multm_compress_rn20;
  assign qs150 = multm_compress_add3b_xor3b_wx149 ^ multm_compress_rn15;
  assign qs151 = multm_compress_add3b_xor3b_wx150 ^ multm_compress_rn5;
  assign qs152 = multm_compress_add3b_xor3b_wx151 ^ multm_compress_rn6;
  assign qs153 = multm_qsp153 ^ multm_qcp152;
  assign qs154 = multm_qsp154 ^ multm_qcp153;
  assign qs155 = multm_compress_add3b_xor3b_wx154 ^ multm_compress_nsd;
  assign qs156 = multm_compress_add3b_xor3b_wx155 ^ multm_compress_ncd;
  assign qs157 = multm_qsp157 ^ multm_qcp156;
  assign qs158 = multm_qsp158 ^ multm_qcp157;
  assign qs159 = multm_qsp159 ^ multm_qcp158;
  assign qs160 = multm_qsp160 ^ multm_qcp159;
  assign qs161 = multm_qsp161 ^ multm_qcp160;
  assign qs162 = multm_compress_add3b_xor3b_wx161 ^ multm_compress_nsd;
  assign qs163 = multm_compress_add3b_xor3b_wx162 ^ multm_compress_ncd;
  assign qs164 = multm_compress_add3b_xor3b_wx163 ^ multm_compress_nsd;
  assign qs165 = multm_compress_add3b_xor3b_wx164 ^ multm_compress_rn4;
  assign qs166 = multm_compress_add3b_xor3b_wx165 ^ multm_compress_rn15;
  assign qs167 = multm_compress_add3b_xor3b_wx166 ^ multm_compress_rn5;
  assign qs168 = multm_compress_add3b_xor3b_wx167 ^ multm_compress_rn20;
  assign qs169 = multm_compress_add3b_xor3b_wx168 ^ multm_compress_rn15;
  assign qs170 = multm_compress_add3b_xor3b_wx169 ^ multm_compress_rn15;
  assign qs171 = multm_compress_add3b_xor3b_wx170 ^ multm_compress_rn15;
  assign qs172 = multm_compress_add3b_xor3b_wx171 ^ multm_compress_rn5;
  assign qs173 = multm_compress_add3b_xor3b_wx172 ^ multm_compress_rn6;
  assign qs174 = multm_qsp174 ^ multm_qcp173;
  assign qs175 = multm_qsp175 ^ multm_qcp174;
  assign qs176 = multm_qsp176 ^ multm_qcp175;
  assign qs177 = multm_compress_add3b_xor3b_wx176 ^ multm_compress_nsd;
  assign qs178 = multm_compress_add3b_xor3b_wx177 ^ multm_compress_rn4;
  assign qs179 = multm_compress_add3b_xor3b_wx178 ^ multm_compress_rn15;
  assign qs180 = multm_compress_add3b_xor3b_wx179 ^ multm_compress_rn5;
  assign qs181 = multm_compress_add3b_xor3b_wx180 ^ multm_compress_rn20;
  assign qs182 = multm_compress_add3b_xor3b_wx181 ^ multm_compress_rn5;
  assign qs183 = multm_compress_add3b_xor3b_wx182 ^ multm_compress_rn6;
  assign san = ~sa;
  assign sap = sb & jp;
  assign saq = san & sap;
  assign sar = ld | saq;
  assign sbp = sa & mdn;
  assign sbq = sb ? jpn : sbp;
  assign sbr = ld | sbq;
  assign srdd = sadd & sbdd;
  assign xn0 = ~multm_jpd;
  assign xn1 = ~multm_reduce_ld1;
  assign xn2 = ~multm_reduce_ld2;
  assign xn3 = ~multm_reduce_pipe0_x5;
  assign xn4 = ~sadd;
  assign xn5 = ~srdd;
  assign xn6 = ~multm_compress_ncd;
  assign dn = dn_o;
  assign ys[0] = ys0_o;
  assign ys[1] = ys1_o;
  assign ys[2] = ys2_o;
  assign ys[3] = ys3_o;
  assign ys[4] = ys4_o;
  assign ys[5] = ys5_o;
  assign ys[6] = ys6_o;
  assign ys[7] = ys7_o;
  assign ys[8] = ys8_o;
  assign ys[9] = ys9_o;
  assign ys[10] = ys10_o;
  assign ys[11] = ys11_o;
  assign ys[12] = ys12_o;
  assign ys[13] = ys13_o;
  assign ys[14] = ys14_o;
  assign ys[15] = ys15_o;
  assign ys[16] = ys16_o;
  assign ys[17] = ys17_o;
  assign ys[18] = ys18_o;
  assign ys[19] = ys19_o;
  assign ys[20] = ys20_o;
  assign ys[21] = ys21_o;
  assign ys[22] = ys22_o;
  assign ys[23] = ys23_o;
  assign ys[24] = ys24_o;
  assign ys[25] = ys25_o;
  assign ys[26] = ys26_o;
  assign ys[27] = ys27_o;
  assign ys[28] = ys28_o;
  assign ys[29] = ys29_o;
  assign ys[30] = ys30_o;
  assign ys[31] = ys31_o;
  assign ys[32] = ys32_o;
  assign ys[33] = ys33_o;
  assign ys[34] = ys34_o;
  assign ys[35] = ys35_o;
  assign ys[36] = ys36_o;
  assign ys[37] = ys37_o;
  assign ys[38] = ys38_o;
  assign ys[39] = ys39_o;
  assign ys[40] = ys40_o;
  assign ys[41] = ys41_o;
  assign ys[42] = ys42_o;
  assign ys[43] = ys43_o;
  assign ys[44] = ys44_o;
  assign ys[45] = ys45_o;
  assign ys[46] = ys46_o;
  assign ys[47] = ys47_o;
  assign ys[48] = ys48_o;
  assign ys[49] = ys49_o;
  assign ys[50] = ys50_o;
  assign ys[51] = ys51_o;
  assign ys[52] = ys52_o;
  assign ys[53] = ys53_o;
  assign ys[54] = ys54_o;
  assign ys[55] = ys55_o;
  assign ys[56] = ys56_o;
  assign ys[57] = ys57_o;
  assign ys[58] = ys58_o;
  assign ys[59] = ys59_o;
  assign ys[60] = ys60_o;
  assign ys[61] = ys61_o;
  assign ys[62] = ys62_o;
  assign ys[63] = ys63_o;
  assign ys[64] = ys64_o;
  assign ys[65] = ys65_o;
  assign ys[66] = ys66_o;
  assign ys[67] = ys67_o;
  assign ys[68] = ys68_o;
  assign ys[69] = ys69_o;
  assign ys[70] = ys70_o;
  assign ys[71] = ys71_o;
  assign ys[72] = ys72_o;
  assign ys[73] = ys73_o;
  assign ys[74] = ys74_o;
  assign ys[75] = ys75_o;
  assign ys[76] = ys76_o;
  assign ys[77] = ys77_o;
  assign ys[78] = ys78_o;
  assign ys[79] = ys79_o;
  assign ys[80] = ys80_o;
  assign ys[81] = ys81_o;
  assign ys[82] = ys82_o;
  assign ys[83] = ys83_o;
  assign ys[84] = ys84_o;
  assign ys[85] = ys85_o;
  assign ys[86] = ys86_o;
  assign ys[87] = ys87_o;
  assign ys[88] = ys88_o;
  assign ys[89] = ys89_o;
  assign ys[90] = ys90_o;
  assign ys[91] = ys91_o;
  assign ys[92] = ys92_o;
  assign ys[93] = ys93_o;
  assign ys[94] = ys94_o;
  assign ys[95] = ys95_o;
  assign ys[96] = ys96_o;
  assign ys[97] = ys97_o;
  assign ys[98] = ys98_o;
  assign ys[99] = ys99_o;
  assign ys[100] = ys100_o;
  assign ys[101] = ys101_o;
  assign ys[102] = ys102_o;
  assign ys[103] = ys103_o;
  assign ys[104] = ys104_o;
  assign ys[105] = ys105_o;
  assign ys[106] = ys106_o;
  assign ys[107] = ys107_o;
  assign ys[108] = ys108_o;
  assign ys[109] = ys109_o;
  assign ys[110] = ys110_o;
  assign ys[111] = ys111_o;
  assign ys[112] = ys112_o;
  assign ys[113] = ys113_o;
  assign ys[114] = ys114_o;
  assign ys[115] = ys115_o;
  assign ys[116] = ys116_o;
  assign ys[117] = ys117_o;
  assign ys[118] = ys118_o;
  assign ys[119] = ys119_o;
  assign ys[120] = ys120_o;
  assign ys[121] = ys121_o;
  assign ys[122] = ys122_o;
  assign ys[123] = ys123_o;
  assign ys[124] = ys124_o;
  assign ys[125] = ys125_o;
  assign ys[126] = ys126_o;
  assign ys[127] = ys127_o;
  assign ys[128] = ys128_o;
  assign ys[129] = ys129_o;
  assign ys[130] = ys130_o;
  assign ys[131] = ys131_o;
  assign ys[132] = ys132_o;
  assign ys[133] = ys133_o;
  assign ys[134] = ys134_o;
  assign ys[135] = ys135_o;
  assign ys[136] = ys136_o;
  assign ys[137] = ys137_o;
  assign ys[138] = ys138_o;
  assign ys[139] = ys139_o;
  assign ys[140] = ys140_o;
  assign ys[141] = ys141_o;
  assign ys[142] = ys142_o;
  assign ys[143] = ys143_o;
  assign ys[144] = ys144_o;
  assign ys[145] = ys145_o;
  assign ys[146] = ys146_o;
  assign ys[147] = ys147_o;
  assign ys[148] = ys148_o;
  assign ys[149] = ys149_o;
  assign ys[150] = ys150_o;
  assign ys[151] = ys151_o;
  assign ys[152] = ys152_o;
  assign ys[153] = ys153_o;
  assign ys[154] = ys154_o;
  assign ys[155] = ys155_o;
  assign ys[156] = ys156_o;
  assign ys[157] = ys157_o;
  assign ys[158] = ys158_o;
  assign ys[159] = ys159_o;
  assign ys[160] = ys160_o;
  assign ys[161] = ys161_o;
  assign ys[162] = ys162_o;
  assign ys[163] = ys163_o;
  assign ys[164] = ys164_o;
  assign ys[165] = ys165_o;
  assign ys[166] = ys166_o;
  assign ys[167] = ys167_o;
  assign ys[168] = ys168_o;
  assign ys[169] = ys169_o;
  assign ys[170] = ys170_o;
  assign ys[171] = ys171_o;
  assign ys[172] = ys172_o;
  assign ys[173] = ys173_o;
  assign ys[174] = ys174_o;
  assign ys[175] = ys175_o;
  assign ys[176] = ys176_o;
  assign ys[177] = ys177_o;
  assign ys[178] = ys178_o;
  assign ys[179] = ys179_o;
  assign ys[180] = ys180_o;
  assign ys[181] = ys181_o;
  assign ys[182] = ys182_o;
  assign ys[183] = ys183_o;
  assign yc[0] = yc0_o;
  assign yc[1] = yc1_o;
  assign yc[2] = yc2_o;
  assign yc[3] = yc3_o;
  assign yc[4] = yc4_o;
  assign yc[5] = yc5_o;
  assign yc[6] = yc6_o;
  assign yc[7] = yc7_o;
  assign yc[8] = yc8_o;
  assign yc[9] = yc9_o;
  assign yc[10] = yc10_o;
  assign yc[11] = yc11_o;
  assign yc[12] = yc12_o;
  assign yc[13] = yc13_o;
  assign yc[14] = yc14_o;
  assign yc[15] = yc15_o;
  assign yc[16] = yc16_o;
  assign yc[17] = yc17_o;
  assign yc[18] = yc18_o;
  assign yc[19] = yc19_o;
  assign yc[20] = yc20_o;
  assign yc[21] = yc21_o;
  assign yc[22] = yc22_o;
  assign yc[23] = yc23_o;
  assign yc[24] = yc24_o;
  assign yc[25] = yc25_o;
  assign yc[26] = yc26_o;
  assign yc[27] = yc27_o;
  assign yc[28] = yc28_o;
  assign yc[29] = yc29_o;
  assign yc[30] = yc30_o;
  assign yc[31] = yc31_o;
  assign yc[32] = yc32_o;
  assign yc[33] = yc33_o;
  assign yc[34] = yc34_o;
  assign yc[35] = yc35_o;
  assign yc[36] = yc36_o;
  assign yc[37] = yc37_o;
  assign yc[38] = yc38_o;
  assign yc[39] = yc39_o;
  assign yc[40] = yc40_o;
  assign yc[41] = yc41_o;
  assign yc[42] = yc42_o;
  assign yc[43] = yc43_o;
  assign yc[44] = yc44_o;
  assign yc[45] = yc45_o;
  assign yc[46] = yc46_o;
  assign yc[47] = yc47_o;
  assign yc[48] = yc48_o;
  assign yc[49] = yc49_o;
  assign yc[50] = yc50_o;
  assign yc[51] = yc51_o;
  assign yc[52] = yc52_o;
  assign yc[53] = yc53_o;
  assign yc[54] = yc54_o;
  assign yc[55] = yc55_o;
  assign yc[56] = yc56_o;
  assign yc[57] = yc57_o;
  assign yc[58] = yc58_o;
  assign yc[59] = yc59_o;
  assign yc[60] = yc60_o;
  assign yc[61] = yc61_o;
  assign yc[62] = yc62_o;
  assign yc[63] = yc63_o;
  assign yc[64] = yc64_o;
  assign yc[65] = yc65_o;
  assign yc[66] = yc66_o;
  assign yc[67] = yc67_o;
  assign yc[68] = yc68_o;
  assign yc[69] = yc69_o;
  assign yc[70] = yc70_o;
  assign yc[71] = yc71_o;
  assign yc[72] = yc72_o;
  assign yc[73] = yc73_o;
  assign yc[74] = yc74_o;
  assign yc[75] = yc75_o;
  assign yc[76] = yc76_o;
  assign yc[77] = yc77_o;
  assign yc[78] = yc78_o;
  assign yc[79] = yc79_o;
  assign yc[80] = yc80_o;
  assign yc[81] = yc81_o;
  assign yc[82] = yc82_o;
  assign yc[83] = yc83_o;
  assign yc[84] = yc84_o;
  assign yc[85] = yc85_o;
  assign yc[86] = yc86_o;
  assign yc[87] = yc87_o;
  assign yc[88] = yc88_o;
  assign yc[89] = yc89_o;
  assign yc[90] = yc90_o;
  assign yc[91] = yc91_o;
  assign yc[92] = yc92_o;
  assign yc[93] = yc93_o;
  assign yc[94] = yc94_o;
  assign yc[95] = yc95_o;
  assign yc[96] = yc96_o;
  assign yc[97] = yc97_o;
  assign yc[98] = yc98_o;
  assign yc[99] = yc99_o;
  assign yc[100] = yc100_o;
  assign yc[101] = yc101_o;
  assign yc[102] = yc102_o;
  assign yc[103] = yc103_o;
  assign yc[104] = yc104_o;
  assign yc[105] = yc105_o;
  assign yc[106] = yc106_o;
  assign yc[107] = yc107_o;
  assign yc[108] = yc108_o;
  assign yc[109] = yc109_o;
  assign yc[110] = yc110_o;
  assign yc[111] = yc111_o;
  assign yc[112] = yc112_o;
  assign yc[113] = yc113_o;
  assign yc[114] = yc114_o;
  assign yc[115] = yc115_o;
  assign yc[116] = yc116_o;
  assign yc[117] = yc117_o;
  assign yc[118] = yc118_o;
  assign yc[119] = yc119_o;
  assign yc[120] = yc120_o;
  assign yc[121] = yc121_o;
  assign yc[122] = yc122_o;
  assign yc[123] = yc123_o;
  assign yc[124] = yc124_o;
  assign yc[125] = yc125_o;
  assign yc[126] = yc126_o;
  assign yc[127] = yc127_o;
  assign yc[128] = yc128_o;
  assign yc[129] = yc129_o;
  assign yc[130] = yc130_o;
  assign yc[131] = yc131_o;
  assign yc[132] = yc132_o;
  assign yc[133] = yc133_o;
  assign yc[134] = yc134_o;
  assign yc[135] = yc135_o;
  assign yc[136] = yc136_o;
  assign yc[137] = yc137_o;
  assign yc[138] = yc138_o;
  assign yc[139] = yc139_o;
  assign yc[140] = yc140_o;
  assign yc[141] = yc141_o;
  assign yc[142] = yc142_o;
  assign yc[143] = yc143_o;
  assign yc[144] = yc144_o;
  assign yc[145] = yc145_o;
  assign yc[146] = yc146_o;
  assign yc[147] = yc147_o;
  assign yc[148] = yc148_o;
  assign yc[149] = yc149_o;
  assign yc[150] = yc150_o;
  assign yc[151] = yc151_o;
  assign yc[152] = yc152_o;
  assign yc[153] = yc153_o;
  assign yc[154] = yc154_o;
  assign yc[155] = yc155_o;
  assign yc[156] = yc156_o;
  assign yc[157] = yc157_o;
  assign yc[158] = yc158_o;
  assign yc[159] = yc159_o;
  assign yc[160] = yc160_o;
  assign yc[161] = yc161_o;
  assign yc[162] = yc162_o;
  assign yc[163] = yc163_o;
  assign yc[164] = yc164_o;
  assign yc[165] = yc165_o;
  assign yc[166] = yc166_o;
  assign yc[167] = yc167_o;
  assign yc[168] = yc168_o;
  assign yc[169] = yc169_o;
  assign yc[170] = yc170_o;
  assign yc[171] = yc171_o;
  assign yc[172] = yc172_o;
  assign yc[173] = yc173_o;
  assign yc[174] = yc174_o;
  assign yc[175] = yc175_o;
  assign yc[176] = yc176_o;
  assign yc[177] = yc177_o;
  assign yc[178] = yc178_o;
  assign yc[179] = yc179_o;
  assign yc[180] = yc180_o;
  assign yc[181] = yc181_o;
  assign yc[182] = yc182_o;
  assign yc[183] = yc183_o;

  always @(posedge clk)
    begin
      ctre_cp0 <= ctre_cr0;
      ctre_cp1 <= ctre_cr1;
      ctre_cp2 <= ctre_cr2;
      ctre_cp3 <= ctre_cr3;
      ctre_cp4 <= ctre_cr4;
      ctre_cp5 <= ctre_cr5;
      ctre_cp6 <= ctre_cr6;
      ctre_cp7 <= ctre_cr7;
      ctre_cp8 <= ctre_cr8;
      ctre_cp9 <= ctre_cr9;
      ctre_dp <= md;
      ctre_sp0 <= ctre_sr0;
      ctre_sp1 <= ctre_sr1;
      ctre_sp2 <= ctre_sr2;
      ctre_sp3 <= ctre_sr3;
      ctre_sp4 <= ctre_sr4;
      ctre_sp5 <= ctre_sr5;
      ctre_sp6 <= ctre_sr6;
      ctre_sp7 <= ctre_sr7;
      ctre_sp8 <= ctre_sr8;
      ctre_sp9 <= ctre_sr9;
      multm_compress_ncd <= multm_compress_pipe1_x4;
      multm_compress_nsd <= multm_compress_pipe0_x4;
      multm_compress_pipe0_x1 <= multm_compress_ns;
      multm_compress_pipe0_x2 <= multm_compress_pipe0_x1;
      multm_compress_pipe0_x3 <= multm_compress_pipe0_x2;
      multm_compress_pipe0_x4 <= multm_compress_pipe0_x3;
      multm_compress_pipe1_x1 <= multm_compress_nc;
      multm_compress_pipe1_x2 <= multm_compress_pipe1_x1;
      multm_compress_pipe1_x3 <= multm_compress_pipe1_x2;
      multm_compress_pipe1_x4 <= multm_compress_pipe1_x3;
      multm_ctrp_ctr_cp0 <= multm_ctrp_ctr_cr0;
      multm_ctrp_ctr_cp1 <= multm_ctrp_ctr_cr1;
      multm_ctrp_ctr_cp2 <= multm_ctrp_ctr_cr2;
      multm_ctrp_ctr_cp3 <= multm_ctrp_ctr_cr3;
      multm_ctrp_ctr_cp4 <= multm_ctrp_ctr_cr4;
      multm_ctrp_ctr_cp5 <= multm_ctrp_ctr_cr5;
      multm_ctrp_ctr_cp6 <= multm_ctrp_ctr_cr6;
      multm_ctrp_ctr_cp7 <= multm_ctrp_ctr_cr7;
      multm_ctrp_ctr_dp <= multm_ctrp_ds;
      multm_ctrp_ctr_sp0 <= multm_ctrp_ctr_sr0;
      multm_ctrp_ctr_sp1 <= multm_ctrp_ctr_sr1;
      multm_ctrp_ctr_sp2 <= multm_ctrp_ctr_sr2;
      multm_ctrp_ctr_sp3 <= multm_ctrp_ctr_sr3;
      multm_ctrp_ctr_sp4 <= multm_ctrp_ctr_sr4;
      multm_ctrp_ctr_sp5 <= multm_ctrp_ctr_sr5;
      multm_ctrp_ctr_sp6 <= multm_ctrp_ctr_sr6;
      multm_jpd <= multm_pipe_x4;
      multm_pipe_x1 <= jp;
      multm_pipe_x2 <= multm_pipe_x1;
      multm_pipe_x3 <= multm_pipe_x2;
      multm_pipe_x4 <= multm_pipe_x3;
      multm_qcp0 <= multm_qcr0;
      multm_qcp1 <= multm_qcr1;
      multm_qcp2 <= multm_qcr2;
      multm_qcp3 <= multm_qcr3;
      multm_qcp4 <= multm_qcr4;
      multm_qcp5 <= multm_qcr5;
      multm_qcp6 <= multm_qcr6;
      multm_qcp7 <= multm_qcr7;
      multm_qcp8 <= multm_qcr8;
      multm_qcp9 <= multm_qcr9;
      multm_qcp10 <= multm_qcr10;
      multm_qcp11 <= multm_qcr11;
      multm_qcp12 <= multm_qcr12;
      multm_qcp13 <= multm_qcr13;
      multm_qcp14 <= multm_qcr14;
      multm_qcp15 <= multm_qcr15;
      multm_qcp16 <= multm_qcr16;
      multm_qcp17 <= multm_qcr17;
      multm_qcp18 <= multm_qcr18;
      multm_qcp19 <= multm_qcr19;
      multm_qcp20 <= multm_qcr20;
      multm_qcp21 <= multm_qcr21;
      multm_qcp22 <= multm_qcr22;
      multm_qcp23 <= multm_qcr23;
      multm_qcp24 <= multm_qcr24;
      multm_qcp25 <= multm_qcr25;
      multm_qcp26 <= multm_qcr26;
      multm_qcp27 <= multm_qcr27;
      multm_qcp28 <= multm_qcr28;
      multm_qcp29 <= multm_qcr29;
      multm_qcp30 <= multm_qcr30;
      multm_qcp31 <= multm_qcr31;
      multm_qcp32 <= multm_qcr32;
      multm_qcp33 <= multm_qcr33;
      multm_qcp34 <= multm_qcr34;
      multm_qcp35 <= multm_qcr35;
      multm_qcp36 <= multm_qcr36;
      multm_qcp37 <= multm_qcr37;
      multm_qcp38 <= multm_qcr38;
      multm_qcp39 <= multm_qcr39;
      multm_qcp40 <= multm_qcr40;
      multm_qcp41 <= multm_qcr41;
      multm_qcp42 <= multm_qcr42;
      multm_qcp43 <= multm_qcr43;
      multm_qcp44 <= multm_qcr44;
      multm_qcp45 <= multm_qcr45;
      multm_qcp46 <= multm_qcr46;
      multm_qcp47 <= multm_qcr47;
      multm_qcp48 <= multm_qcr48;
      multm_qcp49 <= multm_qcr49;
      multm_qcp50 <= multm_qcr50;
      multm_qcp51 <= multm_qcr51;
      multm_qcp52 <= multm_qcr52;
      multm_qcp53 <= multm_qcr53;
      multm_qcp54 <= multm_qcr54;
      multm_qcp55 <= multm_qcr55;
      multm_qcp56 <= multm_qcr56;
      multm_qcp57 <= multm_qcr57;
      multm_qcp58 <= multm_qcr58;
      multm_qcp59 <= multm_qcr59;
      multm_qcp60 <= multm_qcr60;
      multm_qcp61 <= multm_qcr61;
      multm_qcp62 <= multm_qcr62;
      multm_qcp63 <= multm_qcr63;
      multm_qcp64 <= multm_qcr64;
      multm_qcp65 <= multm_qcr65;
      multm_qcp66 <= multm_qcr66;
      multm_qcp67 <= multm_qcr67;
      multm_qcp68 <= multm_qcr68;
      multm_qcp69 <= multm_qcr69;
      multm_qcp70 <= multm_qcr70;
      multm_qcp71 <= multm_qcr71;
      multm_qcp72 <= multm_qcr72;
      multm_qcp73 <= multm_qcr73;
      multm_qcp74 <= multm_qcr74;
      multm_qcp75 <= multm_qcr75;
      multm_qcp76 <= multm_qcr76;
      multm_qcp77 <= multm_qcr77;
      multm_qcp78 <= multm_qcr78;
      multm_qcp79 <= multm_qcr79;
      multm_qcp80 <= multm_qcr80;
      multm_qcp81 <= multm_qcr81;
      multm_qcp82 <= multm_qcr82;
      multm_qcp83 <= multm_qcr83;
      multm_qcp84 <= multm_qcr84;
      multm_qcp85 <= multm_qcr85;
      multm_qcp86 <= multm_qcr86;
      multm_qcp87 <= multm_qcr87;
      multm_qcp88 <= multm_qcr88;
      multm_qcp89 <= multm_qcr89;
      multm_qcp90 <= multm_qcr90;
      multm_qcp91 <= multm_qcr91;
      multm_qcp92 <= multm_qcr92;
      multm_qcp93 <= multm_qcr93;
      multm_qcp94 <= multm_qcr94;
      multm_qcp95 <= multm_qcr95;
      multm_qcp96 <= multm_qcr96;
      multm_qcp97 <= multm_qcr97;
      multm_qcp98 <= multm_qcr98;
      multm_qcp99 <= multm_qcr99;
      multm_qcp100 <= multm_qcr100;
      multm_qcp101 <= multm_qcr101;
      multm_qcp102 <= multm_qcr102;
      multm_qcp103 <= multm_qcr103;
      multm_qcp104 <= multm_qcr104;
      multm_qcp105 <= multm_qcr105;
      multm_qcp106 <= multm_qcr106;
      multm_qcp107 <= multm_qcr107;
      multm_qcp108 <= multm_qcr108;
      multm_qcp109 <= multm_qcr109;
      multm_qcp110 <= multm_qcr110;
      multm_qcp111 <= multm_qcr111;
      multm_qcp112 <= multm_qcr112;
      multm_qcp113 <= multm_qcr113;
      multm_qcp114 <= multm_qcr114;
      multm_qcp115 <= multm_qcr115;
      multm_qcp116 <= multm_qcr116;
      multm_qcp117 <= multm_qcr117;
      multm_qcp118 <= multm_qcr118;
      multm_qcp119 <= multm_qcr119;
      multm_qcp120 <= multm_qcr120;
      multm_qcp121 <= multm_qcr121;
      multm_qcp122 <= multm_qcr122;
      multm_qcp123 <= multm_qcr123;
      multm_qcp124 <= multm_qcr124;
      multm_qcp125 <= multm_qcr125;
      multm_qcp126 <= multm_qcr126;
      multm_qcp127 <= multm_qcr127;
      multm_qcp128 <= multm_qcr128;
      multm_qcp129 <= multm_qcr129;
      multm_qcp130 <= multm_qcr130;
      multm_qcp131 <= multm_qcr131;
      multm_qcp132 <= multm_qcr132;
      multm_qcp133 <= multm_qcr133;
      multm_qcp134 <= multm_qcr134;
      multm_qcp135 <= multm_qcr135;
      multm_qcp136 <= multm_qcr136;
      multm_qcp137 <= multm_qcr137;
      multm_qcp138 <= multm_qcr138;
      multm_qcp139 <= multm_qcr139;
      multm_qcp140 <= multm_qcr140;
      multm_qcp141 <= multm_qcr141;
      multm_qcp142 <= multm_qcr142;
      multm_qcp143 <= multm_qcr143;
      multm_qcp144 <= multm_qcr144;
      multm_qcp145 <= multm_qcr145;
      multm_qcp146 <= multm_qcr146;
      multm_qcp147 <= multm_qcr147;
      multm_qcp148 <= multm_qcr148;
      multm_qcp149 <= multm_qcr149;
      multm_qcp150 <= multm_qcr150;
      multm_qcp151 <= multm_qcr151;
      multm_qcp152 <= multm_qcr152;
      multm_qcp153 <= multm_qcr153;
      multm_qcp154 <= multm_qcr154;
      multm_qcp155 <= multm_qcr155;
      multm_qcp156 <= multm_qcr156;
      multm_qcp157 <= multm_qcr157;
      multm_qcp158 <= multm_qcr158;
      multm_qcp159 <= multm_qcr159;
      multm_qcp160 <= multm_qcr160;
      multm_qcp161 <= multm_qcr161;
      multm_qcp162 <= multm_qcr162;
      multm_qcp163 <= multm_qcr163;
      multm_qcp164 <= multm_qcr164;
      multm_qcp165 <= multm_qcr165;
      multm_qcp166 <= multm_qcr166;
      multm_qcp167 <= multm_qcr167;
      multm_qcp168 <= multm_qcr168;
      multm_qcp169 <= multm_qcr169;
      multm_qcp170 <= multm_qcr170;
      multm_qcp171 <= multm_qcr171;
      multm_qcp172 <= multm_qcr172;
      multm_qcp173 <= multm_qcr173;
      multm_qcp174 <= multm_qcr174;
      multm_qcp175 <= multm_qcr175;
      multm_qcp176 <= multm_qcr176;
      multm_qcp177 <= multm_qcr177;
      multm_qcp178 <= multm_qcr178;
      multm_qcp179 <= multm_qcr179;
      multm_qcp180 <= multm_qcr180;
      multm_qcp181 <= multm_qcr181;
      multm_qcp182 <= multm_qcr182;
      multm_qcp183 <= multm_qcr183;
      multm_qcp184 <= multm_qcr184;
      multm_qsp0 <= multm_qsr0;
      multm_qsp1 <= multm_qsr1;
      multm_qsp2 <= multm_qsr2;
      multm_qsp3 <= multm_qsr3;
      multm_qsp4 <= multm_qsr4;
      multm_qsp5 <= multm_qsr5;
      multm_qsp6 <= multm_qsr6;
      multm_qsp7 <= multm_qsr7;
      multm_qsp8 <= multm_qsr8;
      multm_qsp9 <= multm_qsr9;
      multm_qsp10 <= multm_qsr10;
      multm_qsp11 <= multm_qsr11;
      multm_qsp12 <= multm_qsr12;
      multm_qsp13 <= multm_qsr13;
      multm_qsp14 <= multm_qsr14;
      multm_qsp15 <= multm_qsr15;
      multm_qsp16 <= multm_qsr16;
      multm_qsp17 <= multm_qsr17;
      multm_qsp18 <= multm_qsr18;
      multm_qsp19 <= multm_qsr19;
      multm_qsp20 <= multm_qsr20;
      multm_qsp21 <= multm_qsr21;
      multm_qsp22 <= multm_qsr22;
      multm_qsp23 <= multm_qsr23;
      multm_qsp24 <= multm_qsr24;
      multm_qsp25 <= multm_qsr25;
      multm_qsp26 <= multm_qsr26;
      multm_qsp27 <= multm_qsr27;
      multm_qsp28 <= multm_qsr28;
      multm_qsp29 <= multm_qsr29;
      multm_qsp30 <= multm_qsr30;
      multm_qsp31 <= multm_qsr31;
      multm_qsp32 <= multm_qsr32;
      multm_qsp33 <= multm_qsr33;
      multm_qsp34 <= multm_qsr34;
      multm_qsp35 <= multm_qsr35;
      multm_qsp36 <= multm_qsr36;
      multm_qsp37 <= multm_qsr37;
      multm_qsp38 <= multm_qsr38;
      multm_qsp39 <= multm_qsr39;
      multm_qsp40 <= multm_qsr40;
      multm_qsp41 <= multm_qsr41;
      multm_qsp42 <= multm_qsr42;
      multm_qsp43 <= multm_qsr43;
      multm_qsp44 <= multm_qsr44;
      multm_qsp45 <= multm_qsr45;
      multm_qsp46 <= multm_qsr46;
      multm_qsp47 <= multm_qsr47;
      multm_qsp48 <= multm_qsr48;
      multm_qsp49 <= multm_qsr49;
      multm_qsp50 <= multm_qsr50;
      multm_qsp51 <= multm_qsr51;
      multm_qsp52 <= multm_qsr52;
      multm_qsp53 <= multm_qsr53;
      multm_qsp54 <= multm_qsr54;
      multm_qsp55 <= multm_qsr55;
      multm_qsp56 <= multm_qsr56;
      multm_qsp57 <= multm_qsr57;
      multm_qsp58 <= multm_qsr58;
      multm_qsp59 <= multm_qsr59;
      multm_qsp60 <= multm_qsr60;
      multm_qsp61 <= multm_qsr61;
      multm_qsp62 <= multm_qsr62;
      multm_qsp63 <= multm_qsr63;
      multm_qsp64 <= multm_qsr64;
      multm_qsp65 <= multm_qsr65;
      multm_qsp66 <= multm_qsr66;
      multm_qsp67 <= multm_qsr67;
      multm_qsp68 <= multm_qsr68;
      multm_qsp69 <= multm_qsr69;
      multm_qsp70 <= multm_qsr70;
      multm_qsp71 <= multm_qsr71;
      multm_qsp72 <= multm_qsr72;
      multm_qsp73 <= multm_qsr73;
      multm_qsp74 <= multm_qsr74;
      multm_qsp75 <= multm_qsr75;
      multm_qsp76 <= multm_qsr76;
      multm_qsp77 <= multm_qsr77;
      multm_qsp78 <= multm_qsr78;
      multm_qsp79 <= multm_qsr79;
      multm_qsp80 <= multm_qsr80;
      multm_qsp81 <= multm_qsr81;
      multm_qsp82 <= multm_qsr82;
      multm_qsp83 <= multm_qsr83;
      multm_qsp84 <= multm_qsr84;
      multm_qsp85 <= multm_qsr85;
      multm_qsp86 <= multm_qsr86;
      multm_qsp87 <= multm_qsr87;
      multm_qsp88 <= multm_qsr88;
      multm_qsp89 <= multm_qsr89;
      multm_qsp90 <= multm_qsr90;
      multm_qsp91 <= multm_qsr91;
      multm_qsp92 <= multm_qsr92;
      multm_qsp93 <= multm_qsr93;
      multm_qsp94 <= multm_qsr94;
      multm_qsp95 <= multm_qsr95;
      multm_qsp96 <= multm_qsr96;
      multm_qsp97 <= multm_qsr97;
      multm_qsp98 <= multm_qsr98;
      multm_qsp99 <= multm_qsr99;
      multm_qsp100 <= multm_qsr100;
      multm_qsp101 <= multm_qsr101;
      multm_qsp102 <= multm_qsr102;
      multm_qsp103 <= multm_qsr103;
      multm_qsp104 <= multm_qsr104;
      multm_qsp105 <= multm_qsr105;
      multm_qsp106 <= multm_qsr106;
      multm_qsp107 <= multm_qsr107;
      multm_qsp108 <= multm_qsr108;
      multm_qsp109 <= multm_qsr109;
      multm_qsp110 <= multm_qsr110;
      multm_qsp111 <= multm_qsr111;
      multm_qsp112 <= multm_qsr112;
      multm_qsp113 <= multm_qsr113;
      multm_qsp114 <= multm_qsr114;
      multm_qsp115 <= multm_qsr115;
      multm_qsp116 <= multm_qsr116;
      multm_qsp117 <= multm_qsr117;
      multm_qsp118 <= multm_qsr118;
      multm_qsp119 <= multm_qsr119;
      multm_qsp120 <= multm_qsr120;
      multm_qsp121 <= multm_qsr121;
      multm_qsp122 <= multm_qsr122;
      multm_qsp123 <= multm_qsr123;
      multm_qsp124 <= multm_qsr124;
      multm_qsp125 <= multm_qsr125;
      multm_qsp126 <= multm_qsr126;
      multm_qsp127 <= multm_qsr127;
      multm_qsp128 <= multm_qsr128;
      multm_qsp129 <= multm_qsr129;
      multm_qsp130 <= multm_qsr130;
      multm_qsp131 <= multm_qsr131;
      multm_qsp132 <= multm_qsr132;
      multm_qsp133 <= multm_qsr133;
      multm_qsp134 <= multm_qsr134;
      multm_qsp135 <= multm_qsr135;
      multm_qsp136 <= multm_qsr136;
      multm_qsp137 <= multm_qsr137;
      multm_qsp138 <= multm_qsr138;
      multm_qsp139 <= multm_qsr139;
      multm_qsp140 <= multm_qsr140;
      multm_qsp141 <= multm_qsr141;
      multm_qsp142 <= multm_qsr142;
      multm_qsp143 <= multm_qsr143;
      multm_qsp144 <= multm_qsr144;
      multm_qsp145 <= multm_qsr145;
      multm_qsp146 <= multm_qsr146;
      multm_qsp147 <= multm_qsr147;
      multm_qsp148 <= multm_qsr148;
      multm_qsp149 <= multm_qsr149;
      multm_qsp150 <= multm_qsr150;
      multm_qsp151 <= multm_qsr151;
      multm_qsp152 <= multm_qsr152;
      multm_qsp153 <= multm_qsr153;
      multm_qsp154 <= multm_qsr154;
      multm_qsp155 <= multm_qsr155;
      multm_qsp156 <= multm_qsr156;
      multm_qsp157 <= multm_qsr157;
      multm_qsp158 <= multm_qsr158;
      multm_qsp159 <= multm_qsr159;
      multm_qsp160 <= multm_qsr160;
      multm_qsp161 <= multm_qsr161;
      multm_qsp162 <= multm_qsr162;
      multm_qsp163 <= multm_qsr163;
      multm_qsp164 <= multm_qsr164;
      multm_qsp165 <= multm_qsr165;
      multm_qsp166 <= multm_qsr166;
      multm_qsp167 <= multm_qsr167;
      multm_qsp168 <= multm_qsr168;
      multm_qsp169 <= multm_qsr169;
      multm_qsp170 <= multm_qsr170;
      multm_qsp171 <= multm_qsr171;
      multm_qsp172 <= multm_qsr172;
      multm_qsp173 <= multm_qsr173;
      multm_qsp174 <= multm_qsr174;
      multm_qsp175 <= multm_qsr175;
      multm_qsp176 <= multm_qsr176;
      multm_qsp177 <= multm_qsr177;
      multm_qsp178 <= multm_qsr178;
      multm_qsp179 <= multm_qsr179;
      multm_qsp180 <= multm_qsr180;
      multm_qsp181 <= multm_qsr181;
      multm_qsp182 <= multm_qsr182;
      multm_qsp183 <= multm_qsr183;
      multm_qsp184 <= multm_qsr184;
      multm_reduce_ld1 <= multm_reduce_pipe0_x9;
      multm_reduce_ld2 <= multm_reduce_pipe1_x4;
      multm_reduce_mulb0_cp0 <= multm_reduce_qc0;
      multm_reduce_mulb0_cp1 <= multm_reduce_qc1;
      multm_reduce_mulb0_cp2 <= multm_reduce_qc2;
      multm_reduce_mulb0_cp3 <= multm_reduce_qc3;
      multm_reduce_mulb0_cp4 <= multm_reduce_qc4;
      multm_reduce_mulb0_cp5 <= multm_reduce_qc5;
      multm_reduce_mulb0_cp6 <= multm_reduce_qc6;
      multm_reduce_mulb0_cp7 <= multm_reduce_qc7;
      multm_reduce_mulb0_cp8 <= multm_reduce_qc8;
      multm_reduce_mulb0_cp9 <= multm_reduce_qc9;
      multm_reduce_mulb0_cp10 <= multm_reduce_qc10;
      multm_reduce_mulb0_cp11 <= multm_reduce_qc11;
      multm_reduce_mulb0_cp12 <= multm_reduce_qc12;
      multm_reduce_mulb0_cp13 <= multm_reduce_qc13;
      multm_reduce_mulb0_cp14 <= multm_reduce_qc14;
      multm_reduce_mulb0_cp15 <= multm_reduce_qc15;
      multm_reduce_mulb0_cp16 <= multm_reduce_qc16;
      multm_reduce_mulb0_cp17 <= multm_reduce_qc17;
      multm_reduce_mulb0_cp18 <= multm_reduce_qc18;
      multm_reduce_mulb0_cp19 <= multm_reduce_qc19;
      multm_reduce_mulb0_cp20 <= multm_reduce_qc20;
      multm_reduce_mulb0_cp21 <= multm_reduce_qc21;
      multm_reduce_mulb0_cp22 <= multm_reduce_qc22;
      multm_reduce_mulb0_cp23 <= multm_reduce_qc23;
      multm_reduce_mulb0_cp24 <= multm_reduce_qc24;
      multm_reduce_mulb0_cp25 <= multm_reduce_qc25;
      multm_reduce_mulb0_cp26 <= multm_reduce_qc26;
      multm_reduce_mulb0_cp27 <= multm_reduce_qc27;
      multm_reduce_mulb0_cp28 <= multm_reduce_qc28;
      multm_reduce_mulb0_cp29 <= multm_reduce_qc29;
      multm_reduce_mulb0_cp30 <= multm_reduce_qc30;
      multm_reduce_mulb0_cp31 <= multm_reduce_qc31;
      multm_reduce_mulb0_cp32 <= multm_reduce_qc32;
      multm_reduce_mulb0_cp33 <= multm_reduce_qc33;
      multm_reduce_mulb0_cp34 <= multm_reduce_qc34;
      multm_reduce_mulb0_cp35 <= multm_reduce_qc35;
      multm_reduce_mulb0_cp36 <= multm_reduce_qc36;
      multm_reduce_mulb0_cp37 <= multm_reduce_qc37;
      multm_reduce_mulb0_cp38 <= multm_reduce_qc38;
      multm_reduce_mulb0_cp39 <= multm_reduce_qc39;
      multm_reduce_mulb0_cp40 <= multm_reduce_qc40;
      multm_reduce_mulb0_cp41 <= multm_reduce_qc41;
      multm_reduce_mulb0_cp42 <= multm_reduce_qc42;
      multm_reduce_mulb0_cp43 <= multm_reduce_qc43;
      multm_reduce_mulb0_cp44 <= multm_reduce_qc44;
      multm_reduce_mulb0_cp45 <= multm_reduce_qc45;
      multm_reduce_mulb0_cp46 <= multm_reduce_qc46;
      multm_reduce_mulb0_cp47 <= multm_reduce_qc47;
      multm_reduce_mulb0_cp48 <= multm_reduce_qc48;
      multm_reduce_mulb0_cp49 <= multm_reduce_qc49;
      multm_reduce_mulb0_cp50 <= multm_reduce_qc50;
      multm_reduce_mulb0_cp51 <= multm_reduce_qc51;
      multm_reduce_mulb0_cp52 <= multm_reduce_qc52;
      multm_reduce_mulb0_cp53 <= multm_reduce_qc53;
      multm_reduce_mulb0_cp54 <= multm_reduce_qc54;
      multm_reduce_mulb0_cp55 <= multm_reduce_qc55;
      multm_reduce_mulb0_cp56 <= multm_reduce_qc56;
      multm_reduce_mulb0_cp57 <= multm_reduce_qc57;
      multm_reduce_mulb0_cp58 <= multm_reduce_qc58;
      multm_reduce_mulb0_cp59 <= multm_reduce_qc59;
      multm_reduce_mulb0_cp60 <= multm_reduce_qc60;
      multm_reduce_mulb0_cp61 <= multm_reduce_qc61;
      multm_reduce_mulb0_cp62 <= multm_reduce_qc62;
      multm_reduce_mulb0_cp63 <= multm_reduce_qc63;
      multm_reduce_mulb0_cp64 <= multm_reduce_qc64;
      multm_reduce_mulb0_cp65 <= multm_reduce_qc65;
      multm_reduce_mulb0_cp66 <= multm_reduce_qc66;
      multm_reduce_mulb0_cp67 <= multm_reduce_qc67;
      multm_reduce_mulb0_cp68 <= multm_reduce_qc68;
      multm_reduce_mulb0_cp69 <= multm_reduce_qc69;
      multm_reduce_mulb0_cp70 <= multm_reduce_qc70;
      multm_reduce_mulb0_cp71 <= multm_reduce_qc71;
      multm_reduce_mulb0_cp72 <= multm_reduce_qc72;
      multm_reduce_mulb0_cp73 <= multm_reduce_qc73;
      multm_reduce_mulb0_cp74 <= multm_reduce_qc74;
      multm_reduce_mulb0_cp75 <= multm_reduce_qc75;
      multm_reduce_mulb0_cp76 <= multm_reduce_qc76;
      multm_reduce_mulb0_cp77 <= multm_reduce_qc77;
      multm_reduce_mulb0_cp78 <= multm_reduce_qc78;
      multm_reduce_mulb0_cp79 <= multm_reduce_qc79;
      multm_reduce_mulb0_cp80 <= multm_reduce_qc80;
      multm_reduce_mulb0_cp81 <= multm_reduce_qc81;
      multm_reduce_mulb0_cp82 <= multm_reduce_qc82;
      multm_reduce_mulb0_cp83 <= multm_reduce_qc83;
      multm_reduce_mulb0_cp84 <= multm_reduce_qc84;
      multm_reduce_mulb0_cp85 <= multm_reduce_qc85;
      multm_reduce_mulb0_cp86 <= multm_reduce_qc86;
      multm_reduce_mulb0_cp87 <= multm_reduce_qc87;
      multm_reduce_mulb0_cp88 <= multm_reduce_qc88;
      multm_reduce_mulb0_cp89 <= multm_reduce_qc89;
      multm_reduce_mulb0_cp90 <= multm_reduce_qc90;
      multm_reduce_mulb0_cp91 <= multm_reduce_qc91;
      multm_reduce_mulb0_cp92 <= multm_reduce_qc92;
      multm_reduce_mulb0_cp93 <= multm_reduce_qc93;
      multm_reduce_mulb0_cp94 <= multm_reduce_qc94;
      multm_reduce_mulb0_cp95 <= multm_reduce_qc95;
      multm_reduce_mulb0_cp96 <= multm_reduce_qc96;
      multm_reduce_mulb0_cp97 <= multm_reduce_qc97;
      multm_reduce_mulb0_cp98 <= multm_reduce_qc98;
      multm_reduce_mulb0_cp99 <= multm_reduce_qc99;
      multm_reduce_mulb0_cp100 <= multm_reduce_qc100;
      multm_reduce_mulb0_cp101 <= multm_reduce_qc101;
      multm_reduce_mulb0_cp102 <= multm_reduce_qc102;
      multm_reduce_mulb0_cp103 <= multm_reduce_qc103;
      multm_reduce_mulb0_cp104 <= multm_reduce_qc104;
      multm_reduce_mulb0_cp105 <= multm_reduce_qc105;
      multm_reduce_mulb0_cp106 <= multm_reduce_qc106;
      multm_reduce_mulb0_cp107 <= multm_reduce_qc107;
      multm_reduce_mulb0_cp108 <= multm_reduce_qc108;
      multm_reduce_mulb0_cp109 <= multm_reduce_qc109;
      multm_reduce_mulb0_cp110 <= multm_reduce_qc110;
      multm_reduce_mulb0_cp111 <= multm_reduce_qc111;
      multm_reduce_mulb0_cp112 <= multm_reduce_qc112;
      multm_reduce_mulb0_cp113 <= multm_reduce_qc113;
      multm_reduce_mulb0_cp114 <= multm_reduce_qc114;
      multm_reduce_mulb0_cp115 <= multm_reduce_qc115;
      multm_reduce_mulb0_cp116 <= multm_reduce_qc116;
      multm_reduce_mulb0_cp117 <= multm_reduce_qc117;
      multm_reduce_mulb0_cp118 <= multm_reduce_qc118;
      multm_reduce_mulb0_cp119 <= multm_reduce_qc119;
      multm_reduce_mulb0_cp120 <= multm_reduce_qc120;
      multm_reduce_mulb0_cp121 <= multm_reduce_qc121;
      multm_reduce_mulb0_cp122 <= multm_reduce_qc122;
      multm_reduce_mulb0_cp123 <= multm_reduce_qc123;
      multm_reduce_mulb0_cp124 <= multm_reduce_qc124;
      multm_reduce_mulb0_cp125 <= multm_reduce_qc125;
      multm_reduce_mulb0_cp126 <= multm_reduce_qc126;
      multm_reduce_mulb0_cp127 <= multm_reduce_qc127;
      multm_reduce_mulb0_cp128 <= multm_reduce_qc128;
      multm_reduce_mulb0_cp129 <= multm_reduce_qc129;
      multm_reduce_mulb0_cp130 <= multm_reduce_qc130;
      multm_reduce_mulb0_cp131 <= multm_reduce_qc131;
      multm_reduce_mulb0_cp132 <= multm_reduce_qc132;
      multm_reduce_mulb0_cp133 <= multm_reduce_qc133;
      multm_reduce_mulb0_cp134 <= multm_reduce_qc134;
      multm_reduce_mulb0_cp135 <= multm_reduce_qc135;
      multm_reduce_mulb0_cp136 <= multm_reduce_qc136;
      multm_reduce_mulb0_cp137 <= multm_reduce_qc137;
      multm_reduce_mulb0_cp138 <= multm_reduce_qc138;
      multm_reduce_mulb0_cp139 <= multm_reduce_qc139;
      multm_reduce_mulb0_cp140 <= multm_reduce_qc140;
      multm_reduce_mulb0_cp141 <= multm_reduce_qc141;
      multm_reduce_mulb0_cp142 <= multm_reduce_qc142;
      multm_reduce_mulb0_cp143 <= multm_reduce_qc143;
      multm_reduce_mulb0_cp144 <= multm_reduce_qc144;
      multm_reduce_mulb0_cp145 <= multm_reduce_qc145;
      multm_reduce_mulb0_cp146 <= multm_reduce_qc146;
      multm_reduce_mulb0_cp147 <= multm_reduce_qc147;
      multm_reduce_mulb0_cp148 <= multm_reduce_qc148;
      multm_reduce_mulb0_cp149 <= multm_reduce_qc149;
      multm_reduce_mulb0_cp150 <= multm_reduce_qc150;
      multm_reduce_mulb0_cp151 <= multm_reduce_qc151;
      multm_reduce_mulb0_cp152 <= multm_reduce_qc152;
      multm_reduce_mulb0_cp153 <= multm_reduce_qc153;
      multm_reduce_mulb0_cp154 <= multm_reduce_qc154;
      multm_reduce_mulb0_cp155 <= multm_reduce_qc155;
      multm_reduce_mulb0_cp156 <= multm_reduce_qc156;
      multm_reduce_mulb0_cp157 <= multm_reduce_qc157;
      multm_reduce_mulb0_cp158 <= multm_reduce_qc158;
      multm_reduce_mulb0_cp159 <= multm_reduce_qc159;
      multm_reduce_mulb0_cp160 <= multm_reduce_qc160;
      multm_reduce_mulb0_cp161 <= multm_reduce_qc161;
      multm_reduce_mulb0_cp162 <= multm_reduce_qc162;
      multm_reduce_mulb0_cp163 <= multm_reduce_qc163;
      multm_reduce_mulb0_cp164 <= multm_reduce_qc164;
      multm_reduce_mulb0_cp165 <= multm_reduce_qc165;
      multm_reduce_mulb0_cp166 <= multm_reduce_qc166;
      multm_reduce_mulb0_cp167 <= multm_reduce_qc167;
      multm_reduce_mulb0_cp168 <= multm_reduce_qc168;
      multm_reduce_mulb0_cp169 <= multm_reduce_qc169;
      multm_reduce_mulb0_cp170 <= multm_reduce_qc170;
      multm_reduce_mulb0_cp171 <= multm_reduce_qc171;
      multm_reduce_mulb0_cp172 <= multm_reduce_qc172;
      multm_reduce_mulb0_cp173 <= multm_reduce_qc173;
      multm_reduce_mulb0_cp174 <= multm_reduce_qc174;
      multm_reduce_mulb0_cp175 <= multm_reduce_qc175;
      multm_reduce_mulb0_cp176 <= multm_reduce_qc176;
      multm_reduce_mulb0_cp177 <= multm_reduce_qc177;
      multm_reduce_mulb0_cp178 <= multm_reduce_qc178;
      multm_reduce_mulb0_cp179 <= multm_reduce_qc179;
      multm_reduce_mulb0_cp180 <= multm_reduce_qc180;
      multm_reduce_mulb0_cp181 <= multm_reduce_qc181;
      multm_reduce_mulb0_cp182 <= multm_reduce_qc182;
      multm_reduce_mulb0_cp183 <= multm_reduce_qc183;
      multm_reduce_mulb0_cp184 <= multm_reduce_qc184;
      multm_reduce_mulb0_sp0 <= multm_reduce_qs0;
      multm_reduce_mulb0_sp1 <= multm_reduce_qs1;
      multm_reduce_mulb0_sp2 <= multm_reduce_qs2;
      multm_reduce_mulb0_sp3 <= multm_reduce_qs3;
      multm_reduce_mulb0_sp4 <= multm_reduce_qs4;
      multm_reduce_mulb0_sp5 <= multm_reduce_qs5;
      multm_reduce_mulb0_sp6 <= multm_reduce_qs6;
      multm_reduce_mulb0_sp7 <= multm_reduce_qs7;
      multm_reduce_mulb0_sp8 <= multm_reduce_qs8;
      multm_reduce_mulb0_sp9 <= multm_reduce_qs9;
      multm_reduce_mulb0_sp10 <= multm_reduce_qs10;
      multm_reduce_mulb0_sp11 <= multm_reduce_qs11;
      multm_reduce_mulb0_sp12 <= multm_reduce_qs12;
      multm_reduce_mulb0_sp13 <= multm_reduce_qs13;
      multm_reduce_mulb0_sp14 <= multm_reduce_qs14;
      multm_reduce_mulb0_sp15 <= multm_reduce_qs15;
      multm_reduce_mulb0_sp16 <= multm_reduce_qs16;
      multm_reduce_mulb0_sp17 <= multm_reduce_qs17;
      multm_reduce_mulb0_sp18 <= multm_reduce_qs18;
      multm_reduce_mulb0_sp19 <= multm_reduce_qs19;
      multm_reduce_mulb0_sp20 <= multm_reduce_qs20;
      multm_reduce_mulb0_sp21 <= multm_reduce_qs21;
      multm_reduce_mulb0_sp22 <= multm_reduce_qs22;
      multm_reduce_mulb0_sp23 <= multm_reduce_qs23;
      multm_reduce_mulb0_sp24 <= multm_reduce_qs24;
      multm_reduce_mulb0_sp25 <= multm_reduce_qs25;
      multm_reduce_mulb0_sp26 <= multm_reduce_qs26;
      multm_reduce_mulb0_sp27 <= multm_reduce_qs27;
      multm_reduce_mulb0_sp28 <= multm_reduce_qs28;
      multm_reduce_mulb0_sp29 <= multm_reduce_qs29;
      multm_reduce_mulb0_sp30 <= multm_reduce_qs30;
      multm_reduce_mulb0_sp31 <= multm_reduce_qs31;
      multm_reduce_mulb0_sp32 <= multm_reduce_qs32;
      multm_reduce_mulb0_sp33 <= multm_reduce_qs33;
      multm_reduce_mulb0_sp34 <= multm_reduce_qs34;
      multm_reduce_mulb0_sp35 <= multm_reduce_qs35;
      multm_reduce_mulb0_sp36 <= multm_reduce_qs36;
      multm_reduce_mulb0_sp37 <= multm_reduce_qs37;
      multm_reduce_mulb0_sp38 <= multm_reduce_qs38;
      multm_reduce_mulb0_sp39 <= multm_reduce_qs39;
      multm_reduce_mulb0_sp40 <= multm_reduce_qs40;
      multm_reduce_mulb0_sp41 <= multm_reduce_qs41;
      multm_reduce_mulb0_sp42 <= multm_reduce_qs42;
      multm_reduce_mulb0_sp43 <= multm_reduce_qs43;
      multm_reduce_mulb0_sp44 <= multm_reduce_qs44;
      multm_reduce_mulb0_sp45 <= multm_reduce_qs45;
      multm_reduce_mulb0_sp46 <= multm_reduce_qs46;
      multm_reduce_mulb0_sp47 <= multm_reduce_qs47;
      multm_reduce_mulb0_sp48 <= multm_reduce_qs48;
      multm_reduce_mulb0_sp49 <= multm_reduce_qs49;
      multm_reduce_mulb0_sp50 <= multm_reduce_qs50;
      multm_reduce_mulb0_sp51 <= multm_reduce_qs51;
      multm_reduce_mulb0_sp52 <= multm_reduce_qs52;
      multm_reduce_mulb0_sp53 <= multm_reduce_qs53;
      multm_reduce_mulb0_sp54 <= multm_reduce_qs54;
      multm_reduce_mulb0_sp55 <= multm_reduce_qs55;
      multm_reduce_mulb0_sp56 <= multm_reduce_qs56;
      multm_reduce_mulb0_sp57 <= multm_reduce_qs57;
      multm_reduce_mulb0_sp58 <= multm_reduce_qs58;
      multm_reduce_mulb0_sp59 <= multm_reduce_qs59;
      multm_reduce_mulb0_sp60 <= multm_reduce_qs60;
      multm_reduce_mulb0_sp61 <= multm_reduce_qs61;
      multm_reduce_mulb0_sp62 <= multm_reduce_qs62;
      multm_reduce_mulb0_sp63 <= multm_reduce_qs63;
      multm_reduce_mulb0_sp64 <= multm_reduce_qs64;
      multm_reduce_mulb0_sp65 <= multm_reduce_qs65;
      multm_reduce_mulb0_sp66 <= multm_reduce_qs66;
      multm_reduce_mulb0_sp67 <= multm_reduce_qs67;
      multm_reduce_mulb0_sp68 <= multm_reduce_qs68;
      multm_reduce_mulb0_sp69 <= multm_reduce_qs69;
      multm_reduce_mulb0_sp70 <= multm_reduce_qs70;
      multm_reduce_mulb0_sp71 <= multm_reduce_qs71;
      multm_reduce_mulb0_sp72 <= multm_reduce_qs72;
      multm_reduce_mulb0_sp73 <= multm_reduce_qs73;
      multm_reduce_mulb0_sp74 <= multm_reduce_qs74;
      multm_reduce_mulb0_sp75 <= multm_reduce_qs75;
      multm_reduce_mulb0_sp76 <= multm_reduce_qs76;
      multm_reduce_mulb0_sp77 <= multm_reduce_qs77;
      multm_reduce_mulb0_sp78 <= multm_reduce_qs78;
      multm_reduce_mulb0_sp79 <= multm_reduce_qs79;
      multm_reduce_mulb0_sp80 <= multm_reduce_qs80;
      multm_reduce_mulb0_sp81 <= multm_reduce_qs81;
      multm_reduce_mulb0_sp82 <= multm_reduce_qs82;
      multm_reduce_mulb0_sp83 <= multm_reduce_qs83;
      multm_reduce_mulb0_sp84 <= multm_reduce_qs84;
      multm_reduce_mulb0_sp85 <= multm_reduce_qs85;
      multm_reduce_mulb0_sp86 <= multm_reduce_qs86;
      multm_reduce_mulb0_sp87 <= multm_reduce_qs87;
      multm_reduce_mulb0_sp88 <= multm_reduce_qs88;
      multm_reduce_mulb0_sp89 <= multm_reduce_qs89;
      multm_reduce_mulb0_sp90 <= multm_reduce_qs90;
      multm_reduce_mulb0_sp91 <= multm_reduce_qs91;
      multm_reduce_mulb0_sp92 <= multm_reduce_qs92;
      multm_reduce_mulb0_sp93 <= multm_reduce_qs93;
      multm_reduce_mulb0_sp94 <= multm_reduce_qs94;
      multm_reduce_mulb0_sp95 <= multm_reduce_qs95;
      multm_reduce_mulb0_sp96 <= multm_reduce_qs96;
      multm_reduce_mulb0_sp97 <= multm_reduce_qs97;
      multm_reduce_mulb0_sp98 <= multm_reduce_qs98;
      multm_reduce_mulb0_sp99 <= multm_reduce_qs99;
      multm_reduce_mulb0_sp100 <= multm_reduce_qs100;
      multm_reduce_mulb0_sp101 <= multm_reduce_qs101;
      multm_reduce_mulb0_sp102 <= multm_reduce_qs102;
      multm_reduce_mulb0_sp103 <= multm_reduce_qs103;
      multm_reduce_mulb0_sp104 <= multm_reduce_qs104;
      multm_reduce_mulb0_sp105 <= multm_reduce_qs105;
      multm_reduce_mulb0_sp106 <= multm_reduce_qs106;
      multm_reduce_mulb0_sp107 <= multm_reduce_qs107;
      multm_reduce_mulb0_sp108 <= multm_reduce_qs108;
      multm_reduce_mulb0_sp109 <= multm_reduce_qs109;
      multm_reduce_mulb0_sp110 <= multm_reduce_qs110;
      multm_reduce_mulb0_sp111 <= multm_reduce_qs111;
      multm_reduce_mulb0_sp112 <= multm_reduce_qs112;
      multm_reduce_mulb0_sp113 <= multm_reduce_qs113;
      multm_reduce_mulb0_sp114 <= multm_reduce_qs114;
      multm_reduce_mulb0_sp115 <= multm_reduce_qs115;
      multm_reduce_mulb0_sp116 <= multm_reduce_qs116;
      multm_reduce_mulb0_sp117 <= multm_reduce_qs117;
      multm_reduce_mulb0_sp118 <= multm_reduce_qs118;
      multm_reduce_mulb0_sp119 <= multm_reduce_qs119;
      multm_reduce_mulb0_sp120 <= multm_reduce_qs120;
      multm_reduce_mulb0_sp121 <= multm_reduce_qs121;
      multm_reduce_mulb0_sp122 <= multm_reduce_qs122;
      multm_reduce_mulb0_sp123 <= multm_reduce_qs123;
      multm_reduce_mulb0_sp124 <= multm_reduce_qs124;
      multm_reduce_mulb0_sp125 <= multm_reduce_qs125;
      multm_reduce_mulb0_sp126 <= multm_reduce_qs126;
      multm_reduce_mulb0_sp127 <= multm_reduce_qs127;
      multm_reduce_mulb0_sp128 <= multm_reduce_qs128;
      multm_reduce_mulb0_sp129 <= multm_reduce_qs129;
      multm_reduce_mulb0_sp130 <= multm_reduce_qs130;
      multm_reduce_mulb0_sp131 <= multm_reduce_qs131;
      multm_reduce_mulb0_sp132 <= multm_reduce_qs132;
      multm_reduce_mulb0_sp133 <= multm_reduce_qs133;
      multm_reduce_mulb0_sp134 <= multm_reduce_qs134;
      multm_reduce_mulb0_sp135 <= multm_reduce_qs135;
      multm_reduce_mulb0_sp136 <= multm_reduce_qs136;
      multm_reduce_mulb0_sp137 <= multm_reduce_qs137;
      multm_reduce_mulb0_sp138 <= multm_reduce_qs138;
      multm_reduce_mulb0_sp139 <= multm_reduce_qs139;
      multm_reduce_mulb0_sp140 <= multm_reduce_qs140;
      multm_reduce_mulb0_sp141 <= multm_reduce_qs141;
      multm_reduce_mulb0_sp142 <= multm_reduce_qs142;
      multm_reduce_mulb0_sp143 <= multm_reduce_qs143;
      multm_reduce_mulb0_sp144 <= multm_reduce_qs144;
      multm_reduce_mulb0_sp145 <= multm_reduce_qs145;
      multm_reduce_mulb0_sp146 <= multm_reduce_qs146;
      multm_reduce_mulb0_sp147 <= multm_reduce_qs147;
      multm_reduce_mulb0_sp148 <= multm_reduce_qs148;
      multm_reduce_mulb0_sp149 <= multm_reduce_qs149;
      multm_reduce_mulb0_sp150 <= multm_reduce_qs150;
      multm_reduce_mulb0_sp151 <= multm_reduce_qs151;
      multm_reduce_mulb0_sp152 <= multm_reduce_qs152;
      multm_reduce_mulb0_sp153 <= multm_reduce_qs153;
      multm_reduce_mulb0_sp154 <= multm_reduce_qs154;
      multm_reduce_mulb0_sp155 <= multm_reduce_qs155;
      multm_reduce_mulb0_sp156 <= multm_reduce_qs156;
      multm_reduce_mulb0_sp157 <= multm_reduce_qs157;
      multm_reduce_mulb0_sp158 <= multm_reduce_qs158;
      multm_reduce_mulb0_sp159 <= multm_reduce_qs159;
      multm_reduce_mulb0_sp160 <= multm_reduce_qs160;
      multm_reduce_mulb0_sp161 <= multm_reduce_qs161;
      multm_reduce_mulb0_sp162 <= multm_reduce_qs162;
      multm_reduce_mulb0_sp163 <= multm_reduce_qs163;
      multm_reduce_mulb0_sp164 <= multm_reduce_qs164;
      multm_reduce_mulb0_sp165 <= multm_reduce_qs165;
      multm_reduce_mulb0_sp166 <= multm_reduce_qs166;
      multm_reduce_mulb0_sp167 <= multm_reduce_qs167;
      multm_reduce_mulb0_sp168 <= multm_reduce_qs168;
      multm_reduce_mulb0_sp169 <= multm_reduce_qs169;
      multm_reduce_mulb0_sp170 <= multm_reduce_qs170;
      multm_reduce_mulb0_sp171 <= multm_reduce_qs171;
      multm_reduce_mulb0_sp172 <= multm_reduce_qs172;
      multm_reduce_mulb0_sp173 <= multm_reduce_qs173;
      multm_reduce_mulb0_sp174 <= multm_reduce_qs174;
      multm_reduce_mulb0_sp175 <= multm_reduce_qs175;
      multm_reduce_mulb0_sp176 <= multm_reduce_qs176;
      multm_reduce_mulb0_sp177 <= multm_reduce_qs177;
      multm_reduce_mulb0_sp178 <= multm_reduce_qs178;
      multm_reduce_mulb0_sp179 <= multm_reduce_qs179;
      multm_reduce_mulb0_sp180 <= multm_reduce_qs180;
      multm_reduce_mulb0_sp181 <= multm_reduce_qs181;
      multm_reduce_mulb0_sp182 <= multm_reduce_qs182;
      multm_reduce_mulb0_sp183 <= multm_reduce_qs183;
      multm_reduce_mulb0_sp184 <= multm_reduce_qs184;
      multm_reduce_mulsc_mulb_cp175 <= multm_reduce_pc175;
      multm_reduce_mulsc_mulb_cp176 <= multm_reduce_pc176;
      multm_reduce_mulsc_mulb_cp177 <= multm_reduce_pc177;
      multm_reduce_mulsc_mulb_cp178 <= multm_reduce_pc178;
      multm_reduce_mulsc_mulb_cp179 <= multm_reduce_pc179;
      multm_reduce_mulsc_mulb_cp180 <= multm_reduce_pc180;
      multm_reduce_mulsc_mulb_cp181 <= multm_reduce_pc181;
      multm_reduce_mulsc_mulb_cp182 <= multm_reduce_pc182;
      multm_reduce_mulsc_mulb_cp183 <= multm_reduce_pc183;
      multm_reduce_mulsc_mulb_sp176 <= multm_reduce_ps176;
      multm_reduce_mulsc_mulb_sp177 <= multm_reduce_ps177;
      multm_reduce_mulsc_mulb_sp178 <= multm_reduce_ps178;
      multm_reduce_mulsc_mulb_sp179 <= multm_reduce_ps179;
      multm_reduce_mulsc_mulb_sp180 <= multm_reduce_ps180;
      multm_reduce_mulsc_mulb_sp181 <= multm_reduce_ps181;
      multm_reduce_mulsc_mulb_sp182 <= multm_reduce_ps182;
      multm_reduce_mulsc_mulb_sp183 <= multm_reduce_ps183;
      multm_reduce_mulsc_pipe_x1 <= multm_reduce_mulsc_xb;
      multm_reduce_mulsc_pipe_x2 <= multm_reduce_mulsc_pipe_x1;
      multm_reduce_mulsc_pipe_x3 <= multm_reduce_mulsc_pipe_x2;
      multm_reduce_mulsc_pipe_x4 <= multm_reduce_mulsc_pipe_x3;
      multm_reduce_mulsc_shrsc_cp0 <= multm_reduce_mulsc_shrsc_cr0;
      multm_reduce_mulsc_shrsc_cp1 <= multm_reduce_mulsc_shrsc_cr1;
      multm_reduce_mulsc_shrsc_cp2 <= multm_reduce_mulsc_shrsc_cr2;
      multm_reduce_mulsc_shrsc_cp3 <= multm_reduce_mulsc_shrsc_cr3;
      multm_reduce_mulsc_shrsc_cp4 <= multm_reduce_mulsc_shrsc_cr4;
      multm_reduce_mulsc_shrsc_cp5 <= multm_reduce_mulsc_shrsc_cr5;
      multm_reduce_mulsc_shrsc_cp6 <= multm_reduce_mulsc_shrsc_cr6;
      multm_reduce_mulsc_shrsc_cp7 <= multm_reduce_mulsc_shrsc_cr7;
      multm_reduce_mulsc_shrsc_cp8 <= multm_reduce_mulsc_shrsc_cr8;
      multm_reduce_mulsc_shrsc_cp9 <= multm_reduce_mulsc_shrsc_cr9;
      multm_reduce_mulsc_shrsc_cp10 <= multm_reduce_mulsc_shrsc_cr10;
      multm_reduce_mulsc_shrsc_cp11 <= multm_reduce_mulsc_shrsc_cr11;
      multm_reduce_mulsc_shrsc_cp12 <= multm_reduce_mulsc_shrsc_cr12;
      multm_reduce_mulsc_shrsc_cp13 <= multm_reduce_mulsc_shrsc_cr13;
      multm_reduce_mulsc_shrsc_cp14 <= multm_reduce_mulsc_shrsc_cr14;
      multm_reduce_mulsc_shrsc_cp15 <= multm_reduce_mulsc_shrsc_cr15;
      multm_reduce_mulsc_shrsc_cp16 <= multm_reduce_mulsc_shrsc_cr16;
      multm_reduce_mulsc_shrsc_cp17 <= multm_reduce_mulsc_shrsc_cr17;
      multm_reduce_mulsc_shrsc_cp18 <= multm_reduce_mulsc_shrsc_cr18;
      multm_reduce_mulsc_shrsc_cp19 <= multm_reduce_mulsc_shrsc_cr19;
      multm_reduce_mulsc_shrsc_cp20 <= multm_reduce_mulsc_shrsc_cr20;
      multm_reduce_mulsc_shrsc_cp21 <= multm_reduce_mulsc_shrsc_cr21;
      multm_reduce_mulsc_shrsc_cp22 <= multm_reduce_mulsc_shrsc_cr22;
      multm_reduce_mulsc_shrsc_cp23 <= multm_reduce_mulsc_shrsc_cr23;
      multm_reduce_mulsc_shrsc_cp24 <= multm_reduce_mulsc_shrsc_cr24;
      multm_reduce_mulsc_shrsc_cp25 <= multm_reduce_mulsc_shrsc_cr25;
      multm_reduce_mulsc_shrsc_cp26 <= multm_reduce_mulsc_shrsc_cr26;
      multm_reduce_mulsc_shrsc_cp27 <= multm_reduce_mulsc_shrsc_cr27;
      multm_reduce_mulsc_shrsc_cp28 <= multm_reduce_mulsc_shrsc_cr28;
      multm_reduce_mulsc_shrsc_cp29 <= multm_reduce_mulsc_shrsc_cr29;
      multm_reduce_mulsc_shrsc_cp30 <= multm_reduce_mulsc_shrsc_cr30;
      multm_reduce_mulsc_shrsc_cp31 <= multm_reduce_mulsc_shrsc_cr31;
      multm_reduce_mulsc_shrsc_cp32 <= multm_reduce_mulsc_shrsc_cr32;
      multm_reduce_mulsc_shrsc_cp33 <= multm_reduce_mulsc_shrsc_cr33;
      multm_reduce_mulsc_shrsc_cp34 <= multm_reduce_mulsc_shrsc_cr34;
      multm_reduce_mulsc_shrsc_cp35 <= multm_reduce_mulsc_shrsc_cr35;
      multm_reduce_mulsc_shrsc_cp36 <= multm_reduce_mulsc_shrsc_cr36;
      multm_reduce_mulsc_shrsc_cp37 <= multm_reduce_mulsc_shrsc_cr37;
      multm_reduce_mulsc_shrsc_cp38 <= multm_reduce_mulsc_shrsc_cr38;
      multm_reduce_mulsc_shrsc_cp39 <= multm_reduce_mulsc_shrsc_cr39;
      multm_reduce_mulsc_shrsc_cp40 <= multm_reduce_mulsc_shrsc_cr40;
      multm_reduce_mulsc_shrsc_cp41 <= multm_reduce_mulsc_shrsc_cr41;
      multm_reduce_mulsc_shrsc_cp42 <= multm_reduce_mulsc_shrsc_cr42;
      multm_reduce_mulsc_shrsc_cp43 <= multm_reduce_mulsc_shrsc_cr43;
      multm_reduce_mulsc_shrsc_cp44 <= multm_reduce_mulsc_shrsc_cr44;
      multm_reduce_mulsc_shrsc_cp45 <= multm_reduce_mulsc_shrsc_cr45;
      multm_reduce_mulsc_shrsc_cp46 <= multm_reduce_mulsc_shrsc_cr46;
      multm_reduce_mulsc_shrsc_cp47 <= multm_reduce_mulsc_shrsc_cr47;
      multm_reduce_mulsc_shrsc_cp48 <= multm_reduce_mulsc_shrsc_cr48;
      multm_reduce_mulsc_shrsc_cp49 <= multm_reduce_mulsc_shrsc_cr49;
      multm_reduce_mulsc_shrsc_cp50 <= multm_reduce_mulsc_shrsc_cr50;
      multm_reduce_mulsc_shrsc_cp51 <= multm_reduce_mulsc_shrsc_cr51;
      multm_reduce_mulsc_shrsc_cp52 <= multm_reduce_mulsc_shrsc_cr52;
      multm_reduce_mulsc_shrsc_cp53 <= multm_reduce_mulsc_shrsc_cr53;
      multm_reduce_mulsc_shrsc_cp54 <= multm_reduce_mulsc_shrsc_cr54;
      multm_reduce_mulsc_shrsc_cp55 <= multm_reduce_mulsc_shrsc_cr55;
      multm_reduce_mulsc_shrsc_cp56 <= multm_reduce_mulsc_shrsc_cr56;
      multm_reduce_mulsc_shrsc_cp57 <= multm_reduce_mulsc_shrsc_cr57;
      multm_reduce_mulsc_shrsc_cp58 <= multm_reduce_mulsc_shrsc_cr58;
      multm_reduce_mulsc_shrsc_cp59 <= multm_reduce_mulsc_shrsc_cr59;
      multm_reduce_mulsc_shrsc_cp60 <= multm_reduce_mulsc_shrsc_cr60;
      multm_reduce_mulsc_shrsc_cp61 <= multm_reduce_mulsc_shrsc_cr61;
      multm_reduce_mulsc_shrsc_cp62 <= multm_reduce_mulsc_shrsc_cr62;
      multm_reduce_mulsc_shrsc_cp63 <= multm_reduce_mulsc_shrsc_cr63;
      multm_reduce_mulsc_shrsc_cp64 <= multm_reduce_mulsc_shrsc_cr64;
      multm_reduce_mulsc_shrsc_cp65 <= multm_reduce_mulsc_shrsc_cr65;
      multm_reduce_mulsc_shrsc_cp66 <= multm_reduce_mulsc_shrsc_cr66;
      multm_reduce_mulsc_shrsc_cp67 <= multm_reduce_mulsc_shrsc_cr67;
      multm_reduce_mulsc_shrsc_cp68 <= multm_reduce_mulsc_shrsc_cr68;
      multm_reduce_mulsc_shrsc_cp69 <= multm_reduce_mulsc_shrsc_cr69;
      multm_reduce_mulsc_shrsc_cp70 <= multm_reduce_mulsc_shrsc_cr70;
      multm_reduce_mulsc_shrsc_cp71 <= multm_reduce_mulsc_shrsc_cr71;
      multm_reduce_mulsc_shrsc_cp72 <= multm_reduce_mulsc_shrsc_cr72;
      multm_reduce_mulsc_shrsc_cp73 <= multm_reduce_mulsc_shrsc_cr73;
      multm_reduce_mulsc_shrsc_cp74 <= multm_reduce_mulsc_shrsc_cr74;
      multm_reduce_mulsc_shrsc_cp75 <= multm_reduce_mulsc_shrsc_cr75;
      multm_reduce_mulsc_shrsc_cp76 <= multm_reduce_mulsc_shrsc_cr76;
      multm_reduce_mulsc_shrsc_cp77 <= multm_reduce_mulsc_shrsc_cr77;
      multm_reduce_mulsc_shrsc_cp78 <= multm_reduce_mulsc_shrsc_cr78;
      multm_reduce_mulsc_shrsc_cp79 <= multm_reduce_mulsc_shrsc_cr79;
      multm_reduce_mulsc_shrsc_cp80 <= multm_reduce_mulsc_shrsc_cr80;
      multm_reduce_mulsc_shrsc_cp81 <= multm_reduce_mulsc_shrsc_cr81;
      multm_reduce_mulsc_shrsc_cp82 <= multm_reduce_mulsc_shrsc_cr82;
      multm_reduce_mulsc_shrsc_cp83 <= multm_reduce_mulsc_shrsc_cr83;
      multm_reduce_mulsc_shrsc_cp84 <= multm_reduce_mulsc_shrsc_cr84;
      multm_reduce_mulsc_shrsc_cp85 <= multm_reduce_mulsc_shrsc_cr85;
      multm_reduce_mulsc_shrsc_cp86 <= multm_reduce_mulsc_shrsc_cr86;
      multm_reduce_mulsc_shrsc_cp87 <= multm_reduce_mulsc_shrsc_cr87;
      multm_reduce_mulsc_shrsc_cp88 <= multm_reduce_mulsc_shrsc_cr88;
      multm_reduce_mulsc_shrsc_cp89 <= multm_reduce_mulsc_shrsc_cr89;
      multm_reduce_mulsc_shrsc_cp90 <= multm_reduce_mulsc_shrsc_cr90;
      multm_reduce_mulsc_shrsc_cp91 <= multm_reduce_mulsc_shrsc_cr91;
      multm_reduce_mulsc_shrsc_cp92 <= multm_reduce_mulsc_shrsc_cr92;
      multm_reduce_mulsc_shrsc_cp93 <= multm_reduce_mulsc_shrsc_cr93;
      multm_reduce_mulsc_shrsc_cp94 <= multm_reduce_mulsc_shrsc_cr94;
      multm_reduce_mulsc_shrsc_cp95 <= multm_reduce_mulsc_shrsc_cr95;
      multm_reduce_mulsc_shrsc_cp96 <= multm_reduce_mulsc_shrsc_cr96;
      multm_reduce_mulsc_shrsc_cp97 <= multm_reduce_mulsc_shrsc_cr97;
      multm_reduce_mulsc_shrsc_cp98 <= multm_reduce_mulsc_shrsc_cr98;
      multm_reduce_mulsc_shrsc_cp99 <= multm_reduce_mulsc_shrsc_cr99;
      multm_reduce_mulsc_shrsc_cp100 <= multm_reduce_mulsc_shrsc_cr100;
      multm_reduce_mulsc_shrsc_cp101 <= multm_reduce_mulsc_shrsc_cr101;
      multm_reduce_mulsc_shrsc_cp102 <= multm_reduce_mulsc_shrsc_cr102;
      multm_reduce_mulsc_shrsc_cp103 <= multm_reduce_mulsc_shrsc_cr103;
      multm_reduce_mulsc_shrsc_cp104 <= multm_reduce_mulsc_shrsc_cr104;
      multm_reduce_mulsc_shrsc_cp105 <= multm_reduce_mulsc_shrsc_cr105;
      multm_reduce_mulsc_shrsc_cp106 <= multm_reduce_mulsc_shrsc_cr106;
      multm_reduce_mulsc_shrsc_cp107 <= multm_reduce_mulsc_shrsc_cr107;
      multm_reduce_mulsc_shrsc_cp108 <= multm_reduce_mulsc_shrsc_cr108;
      multm_reduce_mulsc_shrsc_cp109 <= multm_reduce_mulsc_shrsc_cr109;
      multm_reduce_mulsc_shrsc_cp110 <= multm_reduce_mulsc_shrsc_cr110;
      multm_reduce_mulsc_shrsc_cp111 <= multm_reduce_mulsc_shrsc_cr111;
      multm_reduce_mulsc_shrsc_cp112 <= multm_reduce_mulsc_shrsc_cr112;
      multm_reduce_mulsc_shrsc_cp113 <= multm_reduce_mulsc_shrsc_cr113;
      multm_reduce_mulsc_shrsc_cp114 <= multm_reduce_mulsc_shrsc_cr114;
      multm_reduce_mulsc_shrsc_cp115 <= multm_reduce_mulsc_shrsc_cr115;
      multm_reduce_mulsc_shrsc_cp116 <= multm_reduce_mulsc_shrsc_cr116;
      multm_reduce_mulsc_shrsc_cp117 <= multm_reduce_mulsc_shrsc_cr117;
      multm_reduce_mulsc_shrsc_cp118 <= multm_reduce_mulsc_shrsc_cr118;
      multm_reduce_mulsc_shrsc_cp119 <= multm_reduce_mulsc_shrsc_cr119;
      multm_reduce_mulsc_shrsc_cp120 <= multm_reduce_mulsc_shrsc_cr120;
      multm_reduce_mulsc_shrsc_cp121 <= multm_reduce_mulsc_shrsc_cr121;
      multm_reduce_mulsc_shrsc_cp122 <= multm_reduce_mulsc_shrsc_cr122;
      multm_reduce_mulsc_shrsc_cp123 <= multm_reduce_mulsc_shrsc_cr123;
      multm_reduce_mulsc_shrsc_cp124 <= multm_reduce_mulsc_shrsc_cr124;
      multm_reduce_mulsc_shrsc_cp125 <= multm_reduce_mulsc_shrsc_cr125;
      multm_reduce_mulsc_shrsc_cp126 <= multm_reduce_mulsc_shrsc_cr126;
      multm_reduce_mulsc_shrsc_cp127 <= multm_reduce_mulsc_shrsc_cr127;
      multm_reduce_mulsc_shrsc_cp128 <= multm_reduce_mulsc_shrsc_cr128;
      multm_reduce_mulsc_shrsc_cp129 <= multm_reduce_mulsc_shrsc_cr129;
      multm_reduce_mulsc_shrsc_cp130 <= multm_reduce_mulsc_shrsc_cr130;
      multm_reduce_mulsc_shrsc_cp131 <= multm_reduce_mulsc_shrsc_cr131;
      multm_reduce_mulsc_shrsc_cp132 <= multm_reduce_mulsc_shrsc_cr132;
      multm_reduce_mulsc_shrsc_cp133 <= multm_reduce_mulsc_shrsc_cr133;
      multm_reduce_mulsc_shrsc_cp134 <= multm_reduce_mulsc_shrsc_cr134;
      multm_reduce_mulsc_shrsc_cp135 <= multm_reduce_mulsc_shrsc_cr135;
      multm_reduce_mulsc_shrsc_cp136 <= multm_reduce_mulsc_shrsc_cr136;
      multm_reduce_mulsc_shrsc_cp137 <= multm_reduce_mulsc_shrsc_cr137;
      multm_reduce_mulsc_shrsc_cp138 <= multm_reduce_mulsc_shrsc_cr138;
      multm_reduce_mulsc_shrsc_cp139 <= multm_reduce_mulsc_shrsc_cr139;
      multm_reduce_mulsc_shrsc_cp140 <= multm_reduce_mulsc_shrsc_cr140;
      multm_reduce_mulsc_shrsc_cp141 <= multm_reduce_mulsc_shrsc_cr141;
      multm_reduce_mulsc_shrsc_cp142 <= multm_reduce_mulsc_shrsc_cr142;
      multm_reduce_mulsc_shrsc_cp143 <= multm_reduce_mulsc_shrsc_cr143;
      multm_reduce_mulsc_shrsc_cp144 <= multm_reduce_mulsc_shrsc_cr144;
      multm_reduce_mulsc_shrsc_cp145 <= multm_reduce_mulsc_shrsc_cr145;
      multm_reduce_mulsc_shrsc_cp146 <= multm_reduce_mulsc_shrsc_cr146;
      multm_reduce_mulsc_shrsc_cp147 <= multm_reduce_mulsc_shrsc_cr147;
      multm_reduce_mulsc_shrsc_cp148 <= multm_reduce_mulsc_shrsc_cr148;
      multm_reduce_mulsc_shrsc_cp149 <= multm_reduce_mulsc_shrsc_cr149;
      multm_reduce_mulsc_shrsc_cp150 <= multm_reduce_mulsc_shrsc_cr150;
      multm_reduce_mulsc_shrsc_cp151 <= multm_reduce_mulsc_shrsc_cr151;
      multm_reduce_mulsc_shrsc_cp152 <= multm_reduce_mulsc_shrsc_cr152;
      multm_reduce_mulsc_shrsc_cp153 <= multm_reduce_mulsc_shrsc_cr153;
      multm_reduce_mulsc_shrsc_cp154 <= multm_reduce_mulsc_shrsc_cr154;
      multm_reduce_mulsc_shrsc_cp155 <= multm_reduce_mulsc_shrsc_cr155;
      multm_reduce_mulsc_shrsc_cp156 <= multm_reduce_mulsc_shrsc_cr156;
      multm_reduce_mulsc_shrsc_cp157 <= multm_reduce_mulsc_shrsc_cr157;
      multm_reduce_mulsc_shrsc_cp158 <= multm_reduce_mulsc_shrsc_cr158;
      multm_reduce_mulsc_shrsc_cp159 <= multm_reduce_mulsc_shrsc_cr159;
      multm_reduce_mulsc_shrsc_cp160 <= multm_reduce_mulsc_shrsc_cr160;
      multm_reduce_mulsc_shrsc_cp161 <= multm_reduce_mulsc_shrsc_cr161;
      multm_reduce_mulsc_shrsc_cp162 <= multm_reduce_mulsc_shrsc_cr162;
      multm_reduce_mulsc_shrsc_cp163 <= multm_reduce_mulsc_shrsc_cr163;
      multm_reduce_mulsc_shrsc_cp164 <= multm_reduce_mulsc_shrsc_cr164;
      multm_reduce_mulsc_shrsc_cp165 <= multm_reduce_mulsc_shrsc_cr165;
      multm_reduce_mulsc_shrsc_cp166 <= multm_reduce_mulsc_shrsc_cr166;
      multm_reduce_mulsc_shrsc_cp167 <= multm_reduce_mulsc_shrsc_cr167;
      multm_reduce_mulsc_shrsc_cp168 <= multm_reduce_mulsc_shrsc_cr168;
      multm_reduce_mulsc_shrsc_cp169 <= multm_reduce_mulsc_shrsc_cr169;
      multm_reduce_mulsc_shrsc_cp170 <= multm_reduce_mulsc_shrsc_cr170;
      multm_reduce_mulsc_shrsc_cp171 <= multm_reduce_mulsc_shrsc_cr171;
      multm_reduce_mulsc_shrsc_cp172 <= multm_reduce_mulsc_shrsc_cr172;
      multm_reduce_mulsc_shrsc_cp173 <= multm_reduce_mulsc_shrsc_cr173;
      multm_reduce_mulsc_shrsc_cp174 <= multm_reduce_mulsc_shrsc_cr174;
      multm_reduce_mulsc_shrsc_cp175 <= multm_reduce_mulsc_shrsc_cr175;
      multm_reduce_mulsc_shrsc_cp176 <= multm_reduce_mulsc_shrsc_cr176;
      multm_reduce_mulsc_shrsc_cp177 <= multm_reduce_mulsc_shrsc_cr177;
      multm_reduce_mulsc_shrsc_cp178 <= multm_reduce_mulsc_shrsc_cr178;
      multm_reduce_mulsc_shrsc_cp179 <= multm_reduce_mulsc_shrsc_cr179;
      multm_reduce_mulsc_shrsc_cp180 <= multm_reduce_mulsc_shrsc_cr180;
      multm_reduce_mulsc_shrsc_cp181 <= multm_reduce_mulsc_shrsc_cr181;
      multm_reduce_mulsc_shrsc_cp182 <= multm_reduce_mulsc_shrsc_cr182;
      multm_reduce_mulsc_shrsc_cp183 <= multm_reduce_mulsc_shrsc_cr183;
      multm_reduce_mulsc_shrsc_sp0 <= multm_reduce_mulsc_shrsc_sr0;
      multm_reduce_mulsc_shrsc_sp1 <= multm_reduce_mulsc_shrsc_sr1;
      multm_reduce_mulsc_shrsc_sp2 <= multm_reduce_mulsc_shrsc_sr2;
      multm_reduce_mulsc_shrsc_sp3 <= multm_reduce_mulsc_shrsc_sr3;
      multm_reduce_mulsc_shrsc_sp4 <= multm_reduce_mulsc_shrsc_sr4;
      multm_reduce_mulsc_shrsc_sp5 <= multm_reduce_mulsc_shrsc_sr5;
      multm_reduce_mulsc_shrsc_sp6 <= multm_reduce_mulsc_shrsc_sr6;
      multm_reduce_mulsc_shrsc_sp7 <= multm_reduce_mulsc_shrsc_sr7;
      multm_reduce_mulsc_shrsc_sp8 <= multm_reduce_mulsc_shrsc_sr8;
      multm_reduce_mulsc_shrsc_sp9 <= multm_reduce_mulsc_shrsc_sr9;
      multm_reduce_mulsc_shrsc_sp10 <= multm_reduce_mulsc_shrsc_sr10;
      multm_reduce_mulsc_shrsc_sp11 <= multm_reduce_mulsc_shrsc_sr11;
      multm_reduce_mulsc_shrsc_sp12 <= multm_reduce_mulsc_shrsc_sr12;
      multm_reduce_mulsc_shrsc_sp13 <= multm_reduce_mulsc_shrsc_sr13;
      multm_reduce_mulsc_shrsc_sp14 <= multm_reduce_mulsc_shrsc_sr14;
      multm_reduce_mulsc_shrsc_sp15 <= multm_reduce_mulsc_shrsc_sr15;
      multm_reduce_mulsc_shrsc_sp16 <= multm_reduce_mulsc_shrsc_sr16;
      multm_reduce_mulsc_shrsc_sp17 <= multm_reduce_mulsc_shrsc_sr17;
      multm_reduce_mulsc_shrsc_sp18 <= multm_reduce_mulsc_shrsc_sr18;
      multm_reduce_mulsc_shrsc_sp19 <= multm_reduce_mulsc_shrsc_sr19;
      multm_reduce_mulsc_shrsc_sp20 <= multm_reduce_mulsc_shrsc_sr20;
      multm_reduce_mulsc_shrsc_sp21 <= multm_reduce_mulsc_shrsc_sr21;
      multm_reduce_mulsc_shrsc_sp22 <= multm_reduce_mulsc_shrsc_sr22;
      multm_reduce_mulsc_shrsc_sp23 <= multm_reduce_mulsc_shrsc_sr23;
      multm_reduce_mulsc_shrsc_sp24 <= multm_reduce_mulsc_shrsc_sr24;
      multm_reduce_mulsc_shrsc_sp25 <= multm_reduce_mulsc_shrsc_sr25;
      multm_reduce_mulsc_shrsc_sp26 <= multm_reduce_mulsc_shrsc_sr26;
      multm_reduce_mulsc_shrsc_sp27 <= multm_reduce_mulsc_shrsc_sr27;
      multm_reduce_mulsc_shrsc_sp28 <= multm_reduce_mulsc_shrsc_sr28;
      multm_reduce_mulsc_shrsc_sp29 <= multm_reduce_mulsc_shrsc_sr29;
      multm_reduce_mulsc_shrsc_sp30 <= multm_reduce_mulsc_shrsc_sr30;
      multm_reduce_mulsc_shrsc_sp31 <= multm_reduce_mulsc_shrsc_sr31;
      multm_reduce_mulsc_shrsc_sp32 <= multm_reduce_mulsc_shrsc_sr32;
      multm_reduce_mulsc_shrsc_sp33 <= multm_reduce_mulsc_shrsc_sr33;
      multm_reduce_mulsc_shrsc_sp34 <= multm_reduce_mulsc_shrsc_sr34;
      multm_reduce_mulsc_shrsc_sp35 <= multm_reduce_mulsc_shrsc_sr35;
      multm_reduce_mulsc_shrsc_sp36 <= multm_reduce_mulsc_shrsc_sr36;
      multm_reduce_mulsc_shrsc_sp37 <= multm_reduce_mulsc_shrsc_sr37;
      multm_reduce_mulsc_shrsc_sp38 <= multm_reduce_mulsc_shrsc_sr38;
      multm_reduce_mulsc_shrsc_sp39 <= multm_reduce_mulsc_shrsc_sr39;
      multm_reduce_mulsc_shrsc_sp40 <= multm_reduce_mulsc_shrsc_sr40;
      multm_reduce_mulsc_shrsc_sp41 <= multm_reduce_mulsc_shrsc_sr41;
      multm_reduce_mulsc_shrsc_sp42 <= multm_reduce_mulsc_shrsc_sr42;
      multm_reduce_mulsc_shrsc_sp43 <= multm_reduce_mulsc_shrsc_sr43;
      multm_reduce_mulsc_shrsc_sp44 <= multm_reduce_mulsc_shrsc_sr44;
      multm_reduce_mulsc_shrsc_sp45 <= multm_reduce_mulsc_shrsc_sr45;
      multm_reduce_mulsc_shrsc_sp46 <= multm_reduce_mulsc_shrsc_sr46;
      multm_reduce_mulsc_shrsc_sp47 <= multm_reduce_mulsc_shrsc_sr47;
      multm_reduce_mulsc_shrsc_sp48 <= multm_reduce_mulsc_shrsc_sr48;
      multm_reduce_mulsc_shrsc_sp49 <= multm_reduce_mulsc_shrsc_sr49;
      multm_reduce_mulsc_shrsc_sp50 <= multm_reduce_mulsc_shrsc_sr50;
      multm_reduce_mulsc_shrsc_sp51 <= multm_reduce_mulsc_shrsc_sr51;
      multm_reduce_mulsc_shrsc_sp52 <= multm_reduce_mulsc_shrsc_sr52;
      multm_reduce_mulsc_shrsc_sp53 <= multm_reduce_mulsc_shrsc_sr53;
      multm_reduce_mulsc_shrsc_sp54 <= multm_reduce_mulsc_shrsc_sr54;
      multm_reduce_mulsc_shrsc_sp55 <= multm_reduce_mulsc_shrsc_sr55;
      multm_reduce_mulsc_shrsc_sp56 <= multm_reduce_mulsc_shrsc_sr56;
      multm_reduce_mulsc_shrsc_sp57 <= multm_reduce_mulsc_shrsc_sr57;
      multm_reduce_mulsc_shrsc_sp58 <= multm_reduce_mulsc_shrsc_sr58;
      multm_reduce_mulsc_shrsc_sp59 <= multm_reduce_mulsc_shrsc_sr59;
      multm_reduce_mulsc_shrsc_sp60 <= multm_reduce_mulsc_shrsc_sr60;
      multm_reduce_mulsc_shrsc_sp61 <= multm_reduce_mulsc_shrsc_sr61;
      multm_reduce_mulsc_shrsc_sp62 <= multm_reduce_mulsc_shrsc_sr62;
      multm_reduce_mulsc_shrsc_sp63 <= multm_reduce_mulsc_shrsc_sr63;
      multm_reduce_mulsc_shrsc_sp64 <= multm_reduce_mulsc_shrsc_sr64;
      multm_reduce_mulsc_shrsc_sp65 <= multm_reduce_mulsc_shrsc_sr65;
      multm_reduce_mulsc_shrsc_sp66 <= multm_reduce_mulsc_shrsc_sr66;
      multm_reduce_mulsc_shrsc_sp67 <= multm_reduce_mulsc_shrsc_sr67;
      multm_reduce_mulsc_shrsc_sp68 <= multm_reduce_mulsc_shrsc_sr68;
      multm_reduce_mulsc_shrsc_sp69 <= multm_reduce_mulsc_shrsc_sr69;
      multm_reduce_mulsc_shrsc_sp70 <= multm_reduce_mulsc_shrsc_sr70;
      multm_reduce_mulsc_shrsc_sp71 <= multm_reduce_mulsc_shrsc_sr71;
      multm_reduce_mulsc_shrsc_sp72 <= multm_reduce_mulsc_shrsc_sr72;
      multm_reduce_mulsc_shrsc_sp73 <= multm_reduce_mulsc_shrsc_sr73;
      multm_reduce_mulsc_shrsc_sp74 <= multm_reduce_mulsc_shrsc_sr74;
      multm_reduce_mulsc_shrsc_sp75 <= multm_reduce_mulsc_shrsc_sr75;
      multm_reduce_mulsc_shrsc_sp76 <= multm_reduce_mulsc_shrsc_sr76;
      multm_reduce_mulsc_shrsc_sp77 <= multm_reduce_mulsc_shrsc_sr77;
      multm_reduce_mulsc_shrsc_sp78 <= multm_reduce_mulsc_shrsc_sr78;
      multm_reduce_mulsc_shrsc_sp79 <= multm_reduce_mulsc_shrsc_sr79;
      multm_reduce_mulsc_shrsc_sp80 <= multm_reduce_mulsc_shrsc_sr80;
      multm_reduce_mulsc_shrsc_sp81 <= multm_reduce_mulsc_shrsc_sr81;
      multm_reduce_mulsc_shrsc_sp82 <= multm_reduce_mulsc_shrsc_sr82;
      multm_reduce_mulsc_shrsc_sp83 <= multm_reduce_mulsc_shrsc_sr83;
      multm_reduce_mulsc_shrsc_sp84 <= multm_reduce_mulsc_shrsc_sr84;
      multm_reduce_mulsc_shrsc_sp85 <= multm_reduce_mulsc_shrsc_sr85;
      multm_reduce_mulsc_shrsc_sp86 <= multm_reduce_mulsc_shrsc_sr86;
      multm_reduce_mulsc_shrsc_sp87 <= multm_reduce_mulsc_shrsc_sr87;
      multm_reduce_mulsc_shrsc_sp88 <= multm_reduce_mulsc_shrsc_sr88;
      multm_reduce_mulsc_shrsc_sp89 <= multm_reduce_mulsc_shrsc_sr89;
      multm_reduce_mulsc_shrsc_sp90 <= multm_reduce_mulsc_shrsc_sr90;
      multm_reduce_mulsc_shrsc_sp91 <= multm_reduce_mulsc_shrsc_sr91;
      multm_reduce_mulsc_shrsc_sp92 <= multm_reduce_mulsc_shrsc_sr92;
      multm_reduce_mulsc_shrsc_sp93 <= multm_reduce_mulsc_shrsc_sr93;
      multm_reduce_mulsc_shrsc_sp94 <= multm_reduce_mulsc_shrsc_sr94;
      multm_reduce_mulsc_shrsc_sp95 <= multm_reduce_mulsc_shrsc_sr95;
      multm_reduce_mulsc_shrsc_sp96 <= multm_reduce_mulsc_shrsc_sr96;
      multm_reduce_mulsc_shrsc_sp97 <= multm_reduce_mulsc_shrsc_sr97;
      multm_reduce_mulsc_shrsc_sp98 <= multm_reduce_mulsc_shrsc_sr98;
      multm_reduce_mulsc_shrsc_sp99 <= multm_reduce_mulsc_shrsc_sr99;
      multm_reduce_mulsc_shrsc_sp100 <= multm_reduce_mulsc_shrsc_sr100;
      multm_reduce_mulsc_shrsc_sp101 <= multm_reduce_mulsc_shrsc_sr101;
      multm_reduce_mulsc_shrsc_sp102 <= multm_reduce_mulsc_shrsc_sr102;
      multm_reduce_mulsc_shrsc_sp103 <= multm_reduce_mulsc_shrsc_sr103;
      multm_reduce_mulsc_shrsc_sp104 <= multm_reduce_mulsc_shrsc_sr104;
      multm_reduce_mulsc_shrsc_sp105 <= multm_reduce_mulsc_shrsc_sr105;
      multm_reduce_mulsc_shrsc_sp106 <= multm_reduce_mulsc_shrsc_sr106;
      multm_reduce_mulsc_shrsc_sp107 <= multm_reduce_mulsc_shrsc_sr107;
      multm_reduce_mulsc_shrsc_sp108 <= multm_reduce_mulsc_shrsc_sr108;
      multm_reduce_mulsc_shrsc_sp109 <= multm_reduce_mulsc_shrsc_sr109;
      multm_reduce_mulsc_shrsc_sp110 <= multm_reduce_mulsc_shrsc_sr110;
      multm_reduce_mulsc_shrsc_sp111 <= multm_reduce_mulsc_shrsc_sr111;
      multm_reduce_mulsc_shrsc_sp112 <= multm_reduce_mulsc_shrsc_sr112;
      multm_reduce_mulsc_shrsc_sp113 <= multm_reduce_mulsc_shrsc_sr113;
      multm_reduce_mulsc_shrsc_sp114 <= multm_reduce_mulsc_shrsc_sr114;
      multm_reduce_mulsc_shrsc_sp115 <= multm_reduce_mulsc_shrsc_sr115;
      multm_reduce_mulsc_shrsc_sp116 <= multm_reduce_mulsc_shrsc_sr116;
      multm_reduce_mulsc_shrsc_sp117 <= multm_reduce_mulsc_shrsc_sr117;
      multm_reduce_mulsc_shrsc_sp118 <= multm_reduce_mulsc_shrsc_sr118;
      multm_reduce_mulsc_shrsc_sp119 <= multm_reduce_mulsc_shrsc_sr119;
      multm_reduce_mulsc_shrsc_sp120 <= multm_reduce_mulsc_shrsc_sr120;
      multm_reduce_mulsc_shrsc_sp121 <= multm_reduce_mulsc_shrsc_sr121;
      multm_reduce_mulsc_shrsc_sp122 <= multm_reduce_mulsc_shrsc_sr122;
      multm_reduce_mulsc_shrsc_sp123 <= multm_reduce_mulsc_shrsc_sr123;
      multm_reduce_mulsc_shrsc_sp124 <= multm_reduce_mulsc_shrsc_sr124;
      multm_reduce_mulsc_shrsc_sp125 <= multm_reduce_mulsc_shrsc_sr125;
      multm_reduce_mulsc_shrsc_sp126 <= multm_reduce_mulsc_shrsc_sr126;
      multm_reduce_mulsc_shrsc_sp127 <= multm_reduce_mulsc_shrsc_sr127;
      multm_reduce_mulsc_shrsc_sp128 <= multm_reduce_mulsc_shrsc_sr128;
      multm_reduce_mulsc_shrsc_sp129 <= multm_reduce_mulsc_shrsc_sr129;
      multm_reduce_mulsc_shrsc_sp130 <= multm_reduce_mulsc_shrsc_sr130;
      multm_reduce_mulsc_shrsc_sp131 <= multm_reduce_mulsc_shrsc_sr131;
      multm_reduce_mulsc_shrsc_sp132 <= multm_reduce_mulsc_shrsc_sr132;
      multm_reduce_mulsc_shrsc_sp133 <= multm_reduce_mulsc_shrsc_sr133;
      multm_reduce_mulsc_shrsc_sp134 <= multm_reduce_mulsc_shrsc_sr134;
      multm_reduce_mulsc_shrsc_sp135 <= multm_reduce_mulsc_shrsc_sr135;
      multm_reduce_mulsc_shrsc_sp136 <= multm_reduce_mulsc_shrsc_sr136;
      multm_reduce_mulsc_shrsc_sp137 <= multm_reduce_mulsc_shrsc_sr137;
      multm_reduce_mulsc_shrsc_sp138 <= multm_reduce_mulsc_shrsc_sr138;
      multm_reduce_mulsc_shrsc_sp139 <= multm_reduce_mulsc_shrsc_sr139;
      multm_reduce_mulsc_shrsc_sp140 <= multm_reduce_mulsc_shrsc_sr140;
      multm_reduce_mulsc_shrsc_sp141 <= multm_reduce_mulsc_shrsc_sr141;
      multm_reduce_mulsc_shrsc_sp142 <= multm_reduce_mulsc_shrsc_sr142;
      multm_reduce_mulsc_shrsc_sp143 <= multm_reduce_mulsc_shrsc_sr143;
      multm_reduce_mulsc_shrsc_sp144 <= multm_reduce_mulsc_shrsc_sr144;
      multm_reduce_mulsc_shrsc_sp145 <= multm_reduce_mulsc_shrsc_sr145;
      multm_reduce_mulsc_shrsc_sp146 <= multm_reduce_mulsc_shrsc_sr146;
      multm_reduce_mulsc_shrsc_sp147 <= multm_reduce_mulsc_shrsc_sr147;
      multm_reduce_mulsc_shrsc_sp148 <= multm_reduce_mulsc_shrsc_sr148;
      multm_reduce_mulsc_shrsc_sp149 <= multm_reduce_mulsc_shrsc_sr149;
      multm_reduce_mulsc_shrsc_sp150 <= multm_reduce_mulsc_shrsc_sr150;
      multm_reduce_mulsc_shrsc_sp151 <= multm_reduce_mulsc_shrsc_sr151;
      multm_reduce_mulsc_shrsc_sp152 <= multm_reduce_mulsc_shrsc_sr152;
      multm_reduce_mulsc_shrsc_sp153 <= multm_reduce_mulsc_shrsc_sr153;
      multm_reduce_mulsc_shrsc_sp154 <= multm_reduce_mulsc_shrsc_sr154;
      multm_reduce_mulsc_shrsc_sp155 <= multm_reduce_mulsc_shrsc_sr155;
      multm_reduce_mulsc_shrsc_sp156 <= multm_reduce_mulsc_shrsc_sr156;
      multm_reduce_mulsc_shrsc_sp157 <= multm_reduce_mulsc_shrsc_sr157;
      multm_reduce_mulsc_shrsc_sp158 <= multm_reduce_mulsc_shrsc_sr158;
      multm_reduce_mulsc_shrsc_sp159 <= multm_reduce_mulsc_shrsc_sr159;
      multm_reduce_mulsc_shrsc_sp160 <= multm_reduce_mulsc_shrsc_sr160;
      multm_reduce_mulsc_shrsc_sp161 <= multm_reduce_mulsc_shrsc_sr161;
      multm_reduce_mulsc_shrsc_sp162 <= multm_reduce_mulsc_shrsc_sr162;
      multm_reduce_mulsc_shrsc_sp163 <= multm_reduce_mulsc_shrsc_sr163;
      multm_reduce_mulsc_shrsc_sp164 <= multm_reduce_mulsc_shrsc_sr164;
      multm_reduce_mulsc_shrsc_sp165 <= multm_reduce_mulsc_shrsc_sr165;
      multm_reduce_mulsc_shrsc_sp166 <= multm_reduce_mulsc_shrsc_sr166;
      multm_reduce_mulsc_shrsc_sp167 <= multm_reduce_mulsc_shrsc_sr167;
      multm_reduce_mulsc_shrsc_sp168 <= multm_reduce_mulsc_shrsc_sr168;
      multm_reduce_mulsc_shrsc_sp169 <= multm_reduce_mulsc_shrsc_sr169;
      multm_reduce_mulsc_shrsc_sp170 <= multm_reduce_mulsc_shrsc_sr170;
      multm_reduce_mulsc_shrsc_sp171 <= multm_reduce_mulsc_shrsc_sr171;
      multm_reduce_mulsc_shrsc_sp172 <= multm_reduce_mulsc_shrsc_sr172;
      multm_reduce_mulsc_shrsc_sp173 <= multm_reduce_mulsc_shrsc_sr173;
      multm_reduce_mulsc_shrsc_sp174 <= multm_reduce_mulsc_shrsc_sr174;
      multm_reduce_mulsc_shrsc_sp175 <= multm_reduce_mulsc_shrsc_sr175;
      multm_reduce_mulsc_shrsc_sp176 <= multm_reduce_mulsc_shrsc_sr176;
      multm_reduce_mulsc_shrsc_sp177 <= multm_reduce_mulsc_shrsc_sr177;
      multm_reduce_mulsc_shrsc_sp178 <= multm_reduce_mulsc_shrsc_sr178;
      multm_reduce_mulsc_shrsc_sp179 <= multm_reduce_mulsc_shrsc_sr179;
      multm_reduce_mulsc_shrsc_sp180 <= multm_reduce_mulsc_shrsc_sr180;
      multm_reduce_mulsc_shrsc_sp181 <= multm_reduce_mulsc_shrsc_sr181;
      multm_reduce_mulsc_shrsc_sp182 <= multm_reduce_mulsc_shrsc_sr182;
      multm_reduce_mulsc_xbd <= multm_reduce_mulsc_pipe_x4;
      multm_reduce_pipe0_x1 <= sadd;
      multm_reduce_pipe0_x2 <= multm_reduce_pipe0_x1;
      multm_reduce_pipe0_x3 <= multm_reduce_pipe0_x2;
      multm_reduce_pipe0_x4 <= multm_reduce_pipe0_x3;
      multm_reduce_pipe0_x5 <= multm_reduce_pipe0_x4;
      multm_reduce_pipe0_x6 <= multm_reduce_pipe0_x5;
      multm_reduce_pipe0_x7 <= multm_reduce_pipe0_x6;
      multm_reduce_pipe0_x8 <= multm_reduce_pipe0_x7;
      multm_reduce_pipe0_x9 <= multm_reduce_pipe0_x8;
      multm_reduce_pipe1_x1 <= multm_reduce_ld1;
      multm_reduce_pipe1_x2 <= multm_reduce_pipe1_x1;
      multm_reduce_pipe1_x3 <= multm_reduce_pipe1_x2;
      multm_reduce_pipe1_x4 <= multm_reduce_pipe1_x3;
      multm_reduce_pipe2_x1 <= multm_reduce_qb;
      multm_reduce_pipe2_x2 <= multm_reduce_pipe2_x1;
      multm_reduce_pipe2_x3 <= multm_reduce_pipe2_x2;
      multm_reduce_pipe2_x4 <= multm_reduce_pipe2_x3;
      multm_reduce_qb2 <= multm_reduce_pipe2_x4;
      multm_reduce_sa0 <= multm_reduce_sa1;
      multm_reduce_sa1 <= multm_reduce_sa2;
      multm_reduce_sa2 <= multm_reduce_sa3;
      multm_reduce_sa3 <= multm_reduce_sa4;
      multm_reduce_sa4 <= multm_reduce_sa5;
      multm_reduce_sa5 <= multm_reduce_sa6;
      multm_reduce_sa6 <= multm_reduce_sa7;
      multm_reduce_sa7 <= multm_reduce_sa8;
      multm_reduce_sa8 <= multm_reduce_sa9;
      multm_reduce_sa9 <= multm_reduce_pb;
      multm_reduce_sa10 <= multm_reduce_ps0;
      multm_reduce_sa11 <= multm_reduce_ps1;
      multm_reduce_sa12 <= multm_reduce_ps2;
      multm_reduce_sa13 <= multm_reduce_ps3;
      multm_reduce_sa14 <= multm_reduce_ps4;
      multm_reduce_sa15 <= multm_reduce_ps5;
      multm_reduce_sa16 <= multm_reduce_ps6;
      multm_reduce_sa17 <= multm_reduce_ps7;
      multm_reduce_sa18 <= multm_reduce_ps8;
      multm_reduce_sa19 <= multm_reduce_ps9;
      multm_reduce_sa20 <= multm_reduce_ps10;
      multm_reduce_sa21 <= multm_reduce_ps11;
      multm_reduce_sa22 <= multm_reduce_ps12;
      multm_reduce_sa23 <= multm_reduce_ps13;
      multm_reduce_sa24 <= multm_reduce_ps14;
      multm_reduce_sa25 <= multm_reduce_ps15;
      multm_reduce_sa26 <= multm_reduce_ps16;
      multm_reduce_sa27 <= multm_reduce_ps17;
      multm_reduce_sa28 <= multm_reduce_ps18;
      multm_reduce_sa29 <= multm_reduce_ps19;
      multm_reduce_sa30 <= multm_reduce_ps20;
      multm_reduce_sa31 <= multm_reduce_ps21;
      multm_reduce_sa32 <= multm_reduce_ps22;
      multm_reduce_sa33 <= multm_reduce_ps23;
      multm_reduce_sa34 <= multm_reduce_ps24;
      multm_reduce_sa35 <= multm_reduce_ps25;
      multm_reduce_sa36 <= multm_reduce_ps26;
      multm_reduce_sa37 <= multm_reduce_ps27;
      multm_reduce_sa38 <= multm_reduce_ps28;
      multm_reduce_sa39 <= multm_reduce_ps29;
      multm_reduce_sa40 <= multm_reduce_ps30;
      multm_reduce_sa41 <= multm_reduce_ps31;
      multm_reduce_sa42 <= multm_reduce_ps32;
      multm_reduce_sa43 <= multm_reduce_ps33;
      multm_reduce_sa44 <= multm_reduce_ps34;
      multm_reduce_sa45 <= multm_reduce_ps35;
      multm_reduce_sa46 <= multm_reduce_ps36;
      multm_reduce_sa47 <= multm_reduce_ps37;
      multm_reduce_sa48 <= multm_reduce_ps38;
      multm_reduce_sa49 <= multm_reduce_ps39;
      multm_reduce_sa50 <= multm_reduce_ps40;
      multm_reduce_sa51 <= multm_reduce_ps41;
      multm_reduce_sa52 <= multm_reduce_ps42;
      multm_reduce_sa53 <= multm_reduce_ps43;
      multm_reduce_sa54 <= multm_reduce_ps44;
      multm_reduce_sa55 <= multm_reduce_ps45;
      multm_reduce_sa56 <= multm_reduce_ps46;
      multm_reduce_sa57 <= multm_reduce_ps47;
      multm_reduce_sa58 <= multm_reduce_ps48;
      multm_reduce_sa59 <= multm_reduce_ps49;
      multm_reduce_sa60 <= multm_reduce_ps50;
      multm_reduce_sa61 <= multm_reduce_ps51;
      multm_reduce_sa62 <= multm_reduce_ps52;
      multm_reduce_sa63 <= multm_reduce_ps53;
      multm_reduce_sa64 <= multm_reduce_ps54;
      multm_reduce_sa65 <= multm_reduce_ps55;
      multm_reduce_sa66 <= multm_reduce_ps56;
      multm_reduce_sa67 <= multm_reduce_ps57;
      multm_reduce_sa68 <= multm_reduce_ps58;
      multm_reduce_sa69 <= multm_reduce_ps59;
      multm_reduce_sa70 <= multm_reduce_ps60;
      multm_reduce_sa71 <= multm_reduce_ps61;
      multm_reduce_sa72 <= multm_reduce_ps62;
      multm_reduce_sa73 <= multm_reduce_ps63;
      multm_reduce_sa74 <= multm_reduce_ps64;
      multm_reduce_sa75 <= multm_reduce_ps65;
      multm_reduce_sa76 <= multm_reduce_ps66;
      multm_reduce_sa77 <= multm_reduce_ps67;
      multm_reduce_sa78 <= multm_reduce_ps68;
      multm_reduce_sa79 <= multm_reduce_ps69;
      multm_reduce_sa80 <= multm_reduce_ps70;
      multm_reduce_sa81 <= multm_reduce_ps71;
      multm_reduce_sa82 <= multm_reduce_ps72;
      multm_reduce_sa83 <= multm_reduce_ps73;
      multm_reduce_sa84 <= multm_reduce_ps74;
      multm_reduce_sa85 <= multm_reduce_ps75;
      multm_reduce_sa86 <= multm_reduce_ps76;
      multm_reduce_sa87 <= multm_reduce_ps77;
      multm_reduce_sa88 <= multm_reduce_ps78;
      multm_reduce_sa89 <= multm_reduce_ps79;
      multm_reduce_sa90 <= multm_reduce_ps80;
      multm_reduce_sa91 <= multm_reduce_ps81;
      multm_reduce_sa92 <= multm_reduce_ps82;
      multm_reduce_sa93 <= multm_reduce_ps83;
      multm_reduce_sa94 <= multm_reduce_ps84;
      multm_reduce_sa95 <= multm_reduce_ps85;
      multm_reduce_sa96 <= multm_reduce_ps86;
      multm_reduce_sa97 <= multm_reduce_ps87;
      multm_reduce_sa98 <= multm_reduce_ps88;
      multm_reduce_sa99 <= multm_reduce_ps89;
      multm_reduce_sa100 <= multm_reduce_ps90;
      multm_reduce_sa101 <= multm_reduce_ps91;
      multm_reduce_sa102 <= multm_reduce_ps92;
      multm_reduce_sa103 <= multm_reduce_ps93;
      multm_reduce_sa104 <= multm_reduce_ps94;
      multm_reduce_sa105 <= multm_reduce_ps95;
      multm_reduce_sa106 <= multm_reduce_ps96;
      multm_reduce_sa107 <= multm_reduce_ps97;
      multm_reduce_sa108 <= multm_reduce_ps98;
      multm_reduce_sa109 <= multm_reduce_ps99;
      multm_reduce_sa110 <= multm_reduce_ps100;
      multm_reduce_sa111 <= multm_reduce_ps101;
      multm_reduce_sa112 <= multm_reduce_ps102;
      multm_reduce_sa113 <= multm_reduce_ps103;
      multm_reduce_sa114 <= multm_reduce_ps104;
      multm_reduce_sa115 <= multm_reduce_ps105;
      multm_reduce_sa116 <= multm_reduce_ps106;
      multm_reduce_sa117 <= multm_reduce_ps107;
      multm_reduce_sa118 <= multm_reduce_ps108;
      multm_reduce_sa119 <= multm_reduce_ps109;
      multm_reduce_sa120 <= multm_reduce_ps110;
      multm_reduce_sa121 <= multm_reduce_ps111;
      multm_reduce_sa122 <= multm_reduce_ps112;
      multm_reduce_sa123 <= multm_reduce_ps113;
      multm_reduce_sa124 <= multm_reduce_ps114;
      multm_reduce_sa125 <= multm_reduce_ps115;
      multm_reduce_sa126 <= multm_reduce_ps116;
      multm_reduce_sa127 <= multm_reduce_ps117;
      multm_reduce_sa128 <= multm_reduce_ps118;
      multm_reduce_sa129 <= multm_reduce_ps119;
      multm_reduce_sa130 <= multm_reduce_ps120;
      multm_reduce_sa131 <= multm_reduce_ps121;
      multm_reduce_sa132 <= multm_reduce_ps122;
      multm_reduce_sa133 <= multm_reduce_ps123;
      multm_reduce_sa134 <= multm_reduce_ps124;
      multm_reduce_sa135 <= multm_reduce_ps125;
      multm_reduce_sa136 <= multm_reduce_ps126;
      multm_reduce_sa137 <= multm_reduce_ps127;
      multm_reduce_sa138 <= multm_reduce_ps128;
      multm_reduce_sa139 <= multm_reduce_ps129;
      multm_reduce_sa140 <= multm_reduce_ps130;
      multm_reduce_sa141 <= multm_reduce_ps131;
      multm_reduce_sa142 <= multm_reduce_ps132;
      multm_reduce_sa143 <= multm_reduce_ps133;
      multm_reduce_sa144 <= multm_reduce_ps134;
      multm_reduce_sa145 <= multm_reduce_ps135;
      multm_reduce_sa146 <= multm_reduce_ps136;
      multm_reduce_sa147 <= multm_reduce_ps137;
      multm_reduce_sa148 <= multm_reduce_ps138;
      multm_reduce_sa149 <= multm_reduce_ps139;
      multm_reduce_sa150 <= multm_reduce_ps140;
      multm_reduce_sa151 <= multm_reduce_ps141;
      multm_reduce_sa152 <= multm_reduce_ps142;
      multm_reduce_sa153 <= multm_reduce_ps143;
      multm_reduce_sa154 <= multm_reduce_ps144;
      multm_reduce_sa155 <= multm_reduce_ps145;
      multm_reduce_sa156 <= multm_reduce_ps146;
      multm_reduce_sa157 <= multm_reduce_ps147;
      multm_reduce_sa158 <= multm_reduce_ps148;
      multm_reduce_sa159 <= multm_reduce_ps149;
      multm_reduce_sa160 <= multm_reduce_ps150;
      multm_reduce_sa161 <= multm_reduce_ps151;
      multm_reduce_sa162 <= multm_reduce_ps152;
      multm_reduce_sa163 <= multm_reduce_ps153;
      multm_reduce_sa164 <= multm_reduce_ps154;
      multm_reduce_sa165 <= multm_reduce_ps155;
      multm_reduce_sa166 <= multm_reduce_ps156;
      multm_reduce_sa167 <= multm_reduce_ps157;
      multm_reduce_sa168 <= multm_reduce_ps158;
      multm_reduce_sa169 <= multm_reduce_ps159;
      multm_reduce_sa170 <= multm_reduce_ps160;
      multm_reduce_sa171 <= multm_reduce_ps161;
      multm_reduce_sa172 <= multm_reduce_ps162;
      multm_reduce_sa173 <= multm_reduce_ps163;
      multm_reduce_sa174 <= multm_reduce_ps164;
      multm_reduce_sa175 <= multm_reduce_ps165;
      multm_reduce_sa176 <= multm_reduce_ps166;
      multm_reduce_sa177 <= multm_reduce_ps167;
      multm_reduce_sa178 <= multm_reduce_ps168;
      multm_reduce_sa179 <= multm_reduce_ps169;
      multm_reduce_sa180 <= multm_reduce_ps170;
      multm_reduce_sa181 <= multm_reduce_ps171;
      multm_reduce_sa182 <= multm_reduce_ps172;
      multm_reduce_sa183 <= multm_reduce_ps173;
      multm_reduce_sa184 <= multm_reduce_ps174;
      multm_reduce_sa185 <= multm_reduce_ps175;
      multm_reduce_sb0 <= multm_reduce_pc0;
      multm_reduce_sb1 <= multm_reduce_pc1;
      multm_reduce_sb2 <= multm_reduce_pc2;
      multm_reduce_sb3 <= multm_reduce_pc3;
      multm_reduce_sb4 <= multm_reduce_pc4;
      multm_reduce_sb5 <= multm_reduce_pc5;
      multm_reduce_sb6 <= multm_reduce_pc6;
      multm_reduce_sb7 <= multm_reduce_pc7;
      multm_reduce_sb8 <= multm_reduce_pc8;
      multm_reduce_sb9 <= multm_reduce_pc9;
      multm_reduce_sb10 <= multm_reduce_pc10;
      multm_reduce_sb11 <= multm_reduce_pc11;
      multm_reduce_sb12 <= multm_reduce_pc12;
      multm_reduce_sb13 <= multm_reduce_pc13;
      multm_reduce_sb14 <= multm_reduce_pc14;
      multm_reduce_sb15 <= multm_reduce_pc15;
      multm_reduce_sb16 <= multm_reduce_pc16;
      multm_reduce_sb17 <= multm_reduce_pc17;
      multm_reduce_sb18 <= multm_reduce_pc18;
      multm_reduce_sb19 <= multm_reduce_pc19;
      multm_reduce_sb20 <= multm_reduce_pc20;
      multm_reduce_sb21 <= multm_reduce_pc21;
      multm_reduce_sb22 <= multm_reduce_pc22;
      multm_reduce_sb23 <= multm_reduce_pc23;
      multm_reduce_sb24 <= multm_reduce_pc24;
      multm_reduce_sb25 <= multm_reduce_pc25;
      multm_reduce_sb26 <= multm_reduce_pc26;
      multm_reduce_sb27 <= multm_reduce_pc27;
      multm_reduce_sb28 <= multm_reduce_pc28;
      multm_reduce_sb29 <= multm_reduce_pc29;
      multm_reduce_sb30 <= multm_reduce_pc30;
      multm_reduce_sb31 <= multm_reduce_pc31;
      multm_reduce_sb32 <= multm_reduce_pc32;
      multm_reduce_sb33 <= multm_reduce_pc33;
      multm_reduce_sb34 <= multm_reduce_pc34;
      multm_reduce_sb35 <= multm_reduce_pc35;
      multm_reduce_sb36 <= multm_reduce_pc36;
      multm_reduce_sb37 <= multm_reduce_pc37;
      multm_reduce_sb38 <= multm_reduce_pc38;
      multm_reduce_sb39 <= multm_reduce_pc39;
      multm_reduce_sb40 <= multm_reduce_pc40;
      multm_reduce_sb41 <= multm_reduce_pc41;
      multm_reduce_sb42 <= multm_reduce_pc42;
      multm_reduce_sb43 <= multm_reduce_pc43;
      multm_reduce_sb44 <= multm_reduce_pc44;
      multm_reduce_sb45 <= multm_reduce_pc45;
      multm_reduce_sb46 <= multm_reduce_pc46;
      multm_reduce_sb47 <= multm_reduce_pc47;
      multm_reduce_sb48 <= multm_reduce_pc48;
      multm_reduce_sb49 <= multm_reduce_pc49;
      multm_reduce_sb50 <= multm_reduce_pc50;
      multm_reduce_sb51 <= multm_reduce_pc51;
      multm_reduce_sb52 <= multm_reduce_pc52;
      multm_reduce_sb53 <= multm_reduce_pc53;
      multm_reduce_sb54 <= multm_reduce_pc54;
      multm_reduce_sb55 <= multm_reduce_pc55;
      multm_reduce_sb56 <= multm_reduce_pc56;
      multm_reduce_sb57 <= multm_reduce_pc57;
      multm_reduce_sb58 <= multm_reduce_pc58;
      multm_reduce_sb59 <= multm_reduce_pc59;
      multm_reduce_sb60 <= multm_reduce_pc60;
      multm_reduce_sb61 <= multm_reduce_pc61;
      multm_reduce_sb62 <= multm_reduce_pc62;
      multm_reduce_sb63 <= multm_reduce_pc63;
      multm_reduce_sb64 <= multm_reduce_pc64;
      multm_reduce_sb65 <= multm_reduce_pc65;
      multm_reduce_sb66 <= multm_reduce_pc66;
      multm_reduce_sb67 <= multm_reduce_pc67;
      multm_reduce_sb68 <= multm_reduce_pc68;
      multm_reduce_sb69 <= multm_reduce_pc69;
      multm_reduce_sb70 <= multm_reduce_pc70;
      multm_reduce_sb71 <= multm_reduce_pc71;
      multm_reduce_sb72 <= multm_reduce_pc72;
      multm_reduce_sb73 <= multm_reduce_pc73;
      multm_reduce_sb74 <= multm_reduce_pc74;
      multm_reduce_sb75 <= multm_reduce_pc75;
      multm_reduce_sb76 <= multm_reduce_pc76;
      multm_reduce_sb77 <= multm_reduce_pc77;
      multm_reduce_sb78 <= multm_reduce_pc78;
      multm_reduce_sb79 <= multm_reduce_pc79;
      multm_reduce_sb80 <= multm_reduce_pc80;
      multm_reduce_sb81 <= multm_reduce_pc81;
      multm_reduce_sb82 <= multm_reduce_pc82;
      multm_reduce_sb83 <= multm_reduce_pc83;
      multm_reduce_sb84 <= multm_reduce_pc84;
      multm_reduce_sb85 <= multm_reduce_pc85;
      multm_reduce_sb86 <= multm_reduce_pc86;
      multm_reduce_sb87 <= multm_reduce_pc87;
      multm_reduce_sb88 <= multm_reduce_pc88;
      multm_reduce_sb89 <= multm_reduce_pc89;
      multm_reduce_sb90 <= multm_reduce_pc90;
      multm_reduce_sb91 <= multm_reduce_pc91;
      multm_reduce_sb92 <= multm_reduce_pc92;
      multm_reduce_sb93 <= multm_reduce_pc93;
      multm_reduce_sb94 <= multm_reduce_pc94;
      multm_reduce_sb95 <= multm_reduce_pc95;
      multm_reduce_sb96 <= multm_reduce_pc96;
      multm_reduce_sb97 <= multm_reduce_pc97;
      multm_reduce_sb98 <= multm_reduce_pc98;
      multm_reduce_sb99 <= multm_reduce_pc99;
      multm_reduce_sb100 <= multm_reduce_pc100;
      multm_reduce_sb101 <= multm_reduce_pc101;
      multm_reduce_sb102 <= multm_reduce_pc102;
      multm_reduce_sb103 <= multm_reduce_pc103;
      multm_reduce_sb104 <= multm_reduce_pc104;
      multm_reduce_sb105 <= multm_reduce_pc105;
      multm_reduce_sb106 <= multm_reduce_pc106;
      multm_reduce_sb107 <= multm_reduce_pc107;
      multm_reduce_sb108 <= multm_reduce_pc108;
      multm_reduce_sb109 <= multm_reduce_pc109;
      multm_reduce_sb110 <= multm_reduce_pc110;
      multm_reduce_sb111 <= multm_reduce_pc111;
      multm_reduce_sb112 <= multm_reduce_pc112;
      multm_reduce_sb113 <= multm_reduce_pc113;
      multm_reduce_sb114 <= multm_reduce_pc114;
      multm_reduce_sb115 <= multm_reduce_pc115;
      multm_reduce_sb116 <= multm_reduce_pc116;
      multm_reduce_sb117 <= multm_reduce_pc117;
      multm_reduce_sb118 <= multm_reduce_pc118;
      multm_reduce_sb119 <= multm_reduce_pc119;
      multm_reduce_sb120 <= multm_reduce_pc120;
      multm_reduce_sb121 <= multm_reduce_pc121;
      multm_reduce_sb122 <= multm_reduce_pc122;
      multm_reduce_sb123 <= multm_reduce_pc123;
      multm_reduce_sb124 <= multm_reduce_pc124;
      multm_reduce_sb125 <= multm_reduce_pc125;
      multm_reduce_sb126 <= multm_reduce_pc126;
      multm_reduce_sb127 <= multm_reduce_pc127;
      multm_reduce_sb128 <= multm_reduce_pc128;
      multm_reduce_sb129 <= multm_reduce_pc129;
      multm_reduce_sb130 <= multm_reduce_pc130;
      multm_reduce_sb131 <= multm_reduce_pc131;
      multm_reduce_sb132 <= multm_reduce_pc132;
      multm_reduce_sb133 <= multm_reduce_pc133;
      multm_reduce_sb134 <= multm_reduce_pc134;
      multm_reduce_sb135 <= multm_reduce_pc135;
      multm_reduce_sb136 <= multm_reduce_pc136;
      multm_reduce_sb137 <= multm_reduce_pc137;
      multm_reduce_sb138 <= multm_reduce_pc138;
      multm_reduce_sb139 <= multm_reduce_pc139;
      multm_reduce_sb140 <= multm_reduce_pc140;
      multm_reduce_sb141 <= multm_reduce_pc141;
      multm_reduce_sb142 <= multm_reduce_pc142;
      multm_reduce_sb143 <= multm_reduce_pc143;
      multm_reduce_sb144 <= multm_reduce_pc144;
      multm_reduce_sb145 <= multm_reduce_pc145;
      multm_reduce_sb146 <= multm_reduce_pc146;
      multm_reduce_sb147 <= multm_reduce_pc147;
      multm_reduce_sb148 <= multm_reduce_pc148;
      multm_reduce_sb149 <= multm_reduce_pc149;
      multm_reduce_sb150 <= multm_reduce_pc150;
      multm_reduce_sb151 <= multm_reduce_pc151;
      multm_reduce_sb152 <= multm_reduce_pc152;
      multm_reduce_sb153 <= multm_reduce_pc153;
      multm_reduce_sb154 <= multm_reduce_pc154;
      multm_reduce_sb155 <= multm_reduce_pc155;
      multm_reduce_sb156 <= multm_reduce_pc156;
      multm_reduce_sb157 <= multm_reduce_pc157;
      multm_reduce_sb158 <= multm_reduce_pc158;
      multm_reduce_sb159 <= multm_reduce_pc159;
      multm_reduce_sb160 <= multm_reduce_pc160;
      multm_reduce_sb161 <= multm_reduce_pc161;
      multm_reduce_sb162 <= multm_reduce_pc162;
      multm_reduce_sb163 <= multm_reduce_pc163;
      multm_reduce_sb164 <= multm_reduce_pc164;
      multm_reduce_sb165 <= multm_reduce_pc165;
      multm_reduce_sb166 <= multm_reduce_pc166;
      multm_reduce_sb167 <= multm_reduce_pc167;
      multm_reduce_sb168 <= multm_reduce_pc168;
      multm_reduce_sb169 <= multm_reduce_pc169;
      multm_reduce_sb170 <= multm_reduce_pc170;
      multm_reduce_sb171 <= multm_reduce_pc171;
      multm_reduce_sb172 <= multm_reduce_pc172;
      multm_reduce_sb173 <= multm_reduce_pc173;
      multm_reduce_sb174 <= multm_reduce_pc174;
      multm_reduce_sc0 <= multm_reduce_vs0;
      multm_reduce_sc1 <= multm_reduce_vs1;
      multm_reduce_sc2 <= multm_reduce_vs2;
      multm_reduce_sc3 <= multm_reduce_vs3;
      multm_reduce_sc4 <= multm_reduce_vs4;
      multm_reduce_sc5 <= multm_reduce_vs5;
      multm_reduce_sc6 <= multm_reduce_vs6;
      multm_reduce_sc7 <= multm_reduce_vs7;
      multm_reduce_sc8 <= multm_reduce_vs8;
      multm_reduce_sc9 <= multm_reduce_vs9;
      multm_reduce_sc10 <= multm_reduce_vs10;
      multm_reduce_sc11 <= multm_reduce_vs11;
      multm_reduce_sc12 <= multm_reduce_vs12;
      multm_reduce_sc13 <= multm_reduce_vs13;
      multm_reduce_sc14 <= multm_reduce_vs14;
      multm_reduce_sc15 <= multm_reduce_vs15;
      multm_reduce_sc16 <= multm_reduce_vs16;
      multm_reduce_sc17 <= multm_reduce_vs17;
      multm_reduce_sc18 <= multm_reduce_vs18;
      multm_reduce_sc19 <= multm_reduce_vs19;
      multm_reduce_sc20 <= multm_reduce_vs20;
      multm_reduce_sc21 <= multm_reduce_vs21;
      multm_reduce_sc22 <= multm_reduce_vs22;
      multm_reduce_sc23 <= multm_reduce_vs23;
      multm_reduce_sc24 <= multm_reduce_vs24;
      multm_reduce_sc25 <= multm_reduce_vs25;
      multm_reduce_sc26 <= multm_reduce_vs26;
      multm_reduce_sc27 <= multm_reduce_vs27;
      multm_reduce_sc28 <= multm_reduce_vs28;
      multm_reduce_sc29 <= multm_reduce_vs29;
      multm_reduce_sc30 <= multm_reduce_vs30;
      multm_reduce_sc31 <= multm_reduce_vs31;
      multm_reduce_sc32 <= multm_reduce_vs32;
      multm_reduce_sc33 <= multm_reduce_vs33;
      multm_reduce_sc34 <= multm_reduce_vs34;
      multm_reduce_sc35 <= multm_reduce_vs35;
      multm_reduce_sc36 <= multm_reduce_vs36;
      multm_reduce_sc37 <= multm_reduce_vs37;
      multm_reduce_sc38 <= multm_reduce_vs38;
      multm_reduce_sc39 <= multm_reduce_vs39;
      multm_reduce_sc40 <= multm_reduce_vs40;
      multm_reduce_sc41 <= multm_reduce_vs41;
      multm_reduce_sc42 <= multm_reduce_vs42;
      multm_reduce_sc43 <= multm_reduce_vs43;
      multm_reduce_sc44 <= multm_reduce_vs44;
      multm_reduce_sc45 <= multm_reduce_vs45;
      multm_reduce_sc46 <= multm_reduce_vs46;
      multm_reduce_sc47 <= multm_reduce_vs47;
      multm_reduce_sc48 <= multm_reduce_vs48;
      multm_reduce_sc49 <= multm_reduce_vs49;
      multm_reduce_sc50 <= multm_reduce_vs50;
      multm_reduce_sc51 <= multm_reduce_vs51;
      multm_reduce_sc52 <= multm_reduce_vs52;
      multm_reduce_sc53 <= multm_reduce_vs53;
      multm_reduce_sc54 <= multm_reduce_vs54;
      multm_reduce_sc55 <= multm_reduce_vs55;
      multm_reduce_sc56 <= multm_reduce_vs56;
      multm_reduce_sc57 <= multm_reduce_vs57;
      multm_reduce_sc58 <= multm_reduce_vs58;
      multm_reduce_sc59 <= multm_reduce_vs59;
      multm_reduce_sc60 <= multm_reduce_vs60;
      multm_reduce_sc61 <= multm_reduce_vs61;
      multm_reduce_sc62 <= multm_reduce_vs62;
      multm_reduce_sc63 <= multm_reduce_vs63;
      multm_reduce_sc64 <= multm_reduce_vs64;
      multm_reduce_sc65 <= multm_reduce_vs65;
      multm_reduce_sc66 <= multm_reduce_vs66;
      multm_reduce_sc67 <= multm_reduce_vs67;
      multm_reduce_sc68 <= multm_reduce_vs68;
      multm_reduce_sc69 <= multm_reduce_vs69;
      multm_reduce_sc70 <= multm_reduce_vs70;
      multm_reduce_sc71 <= multm_reduce_vs71;
      multm_reduce_sc72 <= multm_reduce_vs72;
      multm_reduce_sc73 <= multm_reduce_vs73;
      multm_reduce_sc74 <= multm_reduce_vs74;
      multm_reduce_sc75 <= multm_reduce_vs75;
      multm_reduce_sc76 <= multm_reduce_vs76;
      multm_reduce_sc77 <= multm_reduce_vs77;
      multm_reduce_sc78 <= multm_reduce_vs78;
      multm_reduce_sc79 <= multm_reduce_vs79;
      multm_reduce_sc80 <= multm_reduce_vs80;
      multm_reduce_sc81 <= multm_reduce_vs81;
      multm_reduce_sc82 <= multm_reduce_vs82;
      multm_reduce_sc83 <= multm_reduce_vs83;
      multm_reduce_sc84 <= multm_reduce_vs84;
      multm_reduce_sc85 <= multm_reduce_vs85;
      multm_reduce_sc86 <= multm_reduce_vs86;
      multm_reduce_sc87 <= multm_reduce_vs87;
      multm_reduce_sc88 <= multm_reduce_vs88;
      multm_reduce_sc89 <= multm_reduce_vs89;
      multm_reduce_sc90 <= multm_reduce_vs90;
      multm_reduce_sc91 <= multm_reduce_vs91;
      multm_reduce_sc92 <= multm_reduce_vs92;
      multm_reduce_sc93 <= multm_reduce_vs93;
      multm_reduce_sc94 <= multm_reduce_vs94;
      multm_reduce_sc95 <= multm_reduce_vs95;
      multm_reduce_sc96 <= multm_reduce_vs96;
      multm_reduce_sc97 <= multm_reduce_vs97;
      multm_reduce_sc98 <= multm_reduce_vs98;
      multm_reduce_sc99 <= multm_reduce_vs99;
      multm_reduce_sc100 <= multm_reduce_vs100;
      multm_reduce_sc101 <= multm_reduce_vs101;
      multm_reduce_sc102 <= multm_reduce_vs102;
      multm_reduce_sc103 <= multm_reduce_vs103;
      multm_reduce_sc104 <= multm_reduce_vs104;
      multm_reduce_sc105 <= multm_reduce_vs105;
      multm_reduce_sc106 <= multm_reduce_vs106;
      multm_reduce_sc107 <= multm_reduce_vs107;
      multm_reduce_sc108 <= multm_reduce_vs108;
      multm_reduce_sc109 <= multm_reduce_vs109;
      multm_reduce_sc110 <= multm_reduce_vs110;
      multm_reduce_sc111 <= multm_reduce_vs111;
      multm_reduce_sc112 <= multm_reduce_vs112;
      multm_reduce_sc113 <= multm_reduce_vs113;
      multm_reduce_sc114 <= multm_reduce_vs114;
      multm_reduce_sc115 <= multm_reduce_vs115;
      multm_reduce_sc116 <= multm_reduce_vs116;
      multm_reduce_sc117 <= multm_reduce_vs117;
      multm_reduce_sc118 <= multm_reduce_vs118;
      multm_reduce_sc119 <= multm_reduce_vs119;
      multm_reduce_sc120 <= multm_reduce_vs120;
      multm_reduce_sc121 <= multm_reduce_vs121;
      multm_reduce_sc122 <= multm_reduce_vs122;
      multm_reduce_sc123 <= multm_reduce_vs123;
      multm_reduce_sc124 <= multm_reduce_vs124;
      multm_reduce_sc125 <= multm_reduce_vs125;
      multm_reduce_sc126 <= multm_reduce_vs126;
      multm_reduce_sc127 <= multm_reduce_vs127;
      multm_reduce_sc128 <= multm_reduce_vs128;
      multm_reduce_sc129 <= multm_reduce_vs129;
      multm_reduce_sc130 <= multm_reduce_vs130;
      multm_reduce_sc131 <= multm_reduce_vs131;
      multm_reduce_sc132 <= multm_reduce_vs132;
      multm_reduce_sc133 <= multm_reduce_vs133;
      multm_reduce_sc134 <= multm_reduce_vs134;
      multm_reduce_sc135 <= multm_reduce_vs135;
      multm_reduce_sc136 <= multm_reduce_vs136;
      multm_reduce_sc137 <= multm_reduce_vs137;
      multm_reduce_sc138 <= multm_reduce_vs138;
      multm_reduce_sc139 <= multm_reduce_vs139;
      multm_reduce_sc140 <= multm_reduce_vs140;
      multm_reduce_sc141 <= multm_reduce_vs141;
      multm_reduce_sc142 <= multm_reduce_vs142;
      multm_reduce_sc143 <= multm_reduce_vs143;
      multm_reduce_sc144 <= multm_reduce_vs144;
      multm_reduce_sc145 <= multm_reduce_vs145;
      multm_reduce_sc146 <= multm_reduce_vs146;
      multm_reduce_sc147 <= multm_reduce_vs147;
      multm_reduce_sc148 <= multm_reduce_vs148;
      multm_reduce_sc149 <= multm_reduce_vs149;
      multm_reduce_sc150 <= multm_reduce_vs150;
      multm_reduce_sc151 <= multm_reduce_vs151;
      multm_reduce_sc152 <= multm_reduce_vs152;
      multm_reduce_sc153 <= multm_reduce_vs153;
      multm_reduce_sc154 <= multm_reduce_vs154;
      multm_reduce_sc155 <= multm_reduce_vs155;
      multm_reduce_sc156 <= multm_reduce_vs156;
      multm_reduce_sc157 <= multm_reduce_vs157;
      multm_reduce_sc158 <= multm_reduce_vs158;
      multm_reduce_sc159 <= multm_reduce_vs159;
      multm_reduce_sc160 <= multm_reduce_vs160;
      multm_reduce_sc161 <= multm_reduce_vs161;
      multm_reduce_sc162 <= multm_reduce_vs162;
      multm_reduce_sc163 <= multm_reduce_vs163;
      multm_reduce_sc164 <= multm_reduce_vs164;
      multm_reduce_sc165 <= multm_reduce_vs165;
      multm_reduce_sc166 <= multm_reduce_vs166;
      multm_reduce_sc167 <= multm_reduce_vs167;
      multm_reduce_sc168 <= multm_reduce_vs168;
      multm_reduce_sc169 <= multm_reduce_vs169;
      multm_reduce_sc170 <= multm_reduce_vs170;
      multm_reduce_sc171 <= multm_reduce_vs171;
      multm_reduce_sc172 <= multm_reduce_vs172;
      multm_reduce_sc173 <= multm_reduce_vs173;
      multm_reduce_sc174 <= multm_reduce_vs174;
      multm_reduce_sc175 <= multm_reduce_vs175;
      multm_reduce_sc176 <= multm_reduce_vs176;
      multm_reduce_sc177 <= multm_reduce_vs177;
      multm_reduce_sc178 <= multm_reduce_vs178;
      multm_reduce_sc179 <= multm_reduce_vs179;
      multm_reduce_sc180 <= multm_reduce_vs180;
      multm_reduce_sc181 <= multm_reduce_vs181;
      multm_reduce_sc182 <= multm_reduce_vs182;
      multm_reduce_sd0 <= multm_reduce_vt;
      multm_reduce_sd1 <= multm_reduce_vc0;
      multm_reduce_sd2 <= multm_reduce_vc1;
      multm_reduce_sd3 <= multm_reduce_vc2;
      multm_reduce_sd4 <= multm_reduce_vc3;
      multm_reduce_sd5 <= multm_reduce_vc4;
      multm_reduce_sd6 <= multm_reduce_vc5;
      multm_reduce_sd7 <= multm_reduce_vc6;
      multm_reduce_sd8 <= multm_reduce_vc7;
      multm_reduce_sd9 <= multm_reduce_vc8;
      multm_reduce_sd10 <= multm_reduce_vc9;
      multm_reduce_sd11 <= multm_reduce_vc10;
      multm_reduce_sd12 <= multm_reduce_vc11;
      multm_reduce_sd13 <= multm_reduce_vc12;
      multm_reduce_sd14 <= multm_reduce_vc13;
      multm_reduce_sd15 <= multm_reduce_vc14;
      multm_reduce_sd16 <= multm_reduce_vc15;
      multm_reduce_sd17 <= multm_reduce_vc16;
      multm_reduce_sd18 <= multm_reduce_vc17;
      multm_reduce_sd19 <= multm_reduce_vc18;
      multm_reduce_sd20 <= multm_reduce_vc19;
      multm_reduce_sd21 <= multm_reduce_vc20;
      multm_reduce_sd22 <= multm_reduce_vc21;
      multm_reduce_sd23 <= multm_reduce_vc22;
      multm_reduce_sd24 <= multm_reduce_vc23;
      multm_reduce_sd25 <= multm_reduce_vc24;
      multm_reduce_sd26 <= multm_reduce_vc25;
      multm_reduce_sd27 <= multm_reduce_vc26;
      multm_reduce_sd28 <= multm_reduce_vc27;
      multm_reduce_sd29 <= multm_reduce_vc28;
      multm_reduce_sd30 <= multm_reduce_vc29;
      multm_reduce_sd31 <= multm_reduce_vc30;
      multm_reduce_sd32 <= multm_reduce_vc31;
      multm_reduce_sd33 <= multm_reduce_vc32;
      multm_reduce_sd34 <= multm_reduce_vc33;
      multm_reduce_sd35 <= multm_reduce_vc34;
      multm_reduce_sd36 <= multm_reduce_vc35;
      multm_reduce_sd37 <= multm_reduce_vc36;
      multm_reduce_sd38 <= multm_reduce_vc37;
      multm_reduce_sd39 <= multm_reduce_vc38;
      multm_reduce_sd40 <= multm_reduce_vc39;
      multm_reduce_sd41 <= multm_reduce_vc40;
      multm_reduce_sd42 <= multm_reduce_vc41;
      multm_reduce_sd43 <= multm_reduce_vc42;
      multm_reduce_sd44 <= multm_reduce_vc43;
      multm_reduce_sd45 <= multm_reduce_vc44;
      multm_reduce_sd46 <= multm_reduce_vc45;
      multm_reduce_sd47 <= multm_reduce_vc46;
      multm_reduce_sd48 <= multm_reduce_vc47;
      multm_reduce_sd49 <= multm_reduce_vc48;
      multm_reduce_sd50 <= multm_reduce_vc49;
      multm_reduce_sd51 <= multm_reduce_vc50;
      multm_reduce_sd52 <= multm_reduce_vc51;
      multm_reduce_sd53 <= multm_reduce_vc52;
      multm_reduce_sd54 <= multm_reduce_vc53;
      multm_reduce_sd55 <= multm_reduce_vc54;
      multm_reduce_sd56 <= multm_reduce_vc55;
      multm_reduce_sd57 <= multm_reduce_vc56;
      multm_reduce_sd58 <= multm_reduce_vc57;
      multm_reduce_sd59 <= multm_reduce_vc58;
      multm_reduce_sd60 <= multm_reduce_vc59;
      multm_reduce_sd61 <= multm_reduce_vc60;
      multm_reduce_sd62 <= multm_reduce_vc61;
      multm_reduce_sd63 <= multm_reduce_vc62;
      multm_reduce_sd64 <= multm_reduce_vc63;
      multm_reduce_sd65 <= multm_reduce_vc64;
      multm_reduce_sd66 <= multm_reduce_vc65;
      multm_reduce_sd67 <= multm_reduce_vc66;
      multm_reduce_sd68 <= multm_reduce_vc67;
      multm_reduce_sd69 <= multm_reduce_vc68;
      multm_reduce_sd70 <= multm_reduce_vc69;
      multm_reduce_sd71 <= multm_reduce_vc70;
      multm_reduce_sd72 <= multm_reduce_vc71;
      multm_reduce_sd73 <= multm_reduce_vc72;
      multm_reduce_sd74 <= multm_reduce_vc73;
      multm_reduce_sd75 <= multm_reduce_vc74;
      multm_reduce_sd76 <= multm_reduce_vc75;
      multm_reduce_sd77 <= multm_reduce_vc76;
      multm_reduce_sd78 <= multm_reduce_vc77;
      multm_reduce_sd79 <= multm_reduce_vc78;
      multm_reduce_sd80 <= multm_reduce_vc79;
      multm_reduce_sd81 <= multm_reduce_vc80;
      multm_reduce_sd82 <= multm_reduce_vc81;
      multm_reduce_sd83 <= multm_reduce_vc82;
      multm_reduce_sd84 <= multm_reduce_vc83;
      multm_reduce_sd85 <= multm_reduce_vc84;
      multm_reduce_sd86 <= multm_reduce_vc85;
      multm_reduce_sd87 <= multm_reduce_vc86;
      multm_reduce_sd88 <= multm_reduce_vc87;
      multm_reduce_sd89 <= multm_reduce_vc88;
      multm_reduce_sd90 <= multm_reduce_vc89;
      multm_reduce_sd91 <= multm_reduce_vc90;
      multm_reduce_sd92 <= multm_reduce_vc91;
      multm_reduce_sd93 <= multm_reduce_vc92;
      multm_reduce_sd94 <= multm_reduce_vc93;
      multm_reduce_sd95 <= multm_reduce_vc94;
      multm_reduce_sd96 <= multm_reduce_vc95;
      multm_reduce_sd97 <= multm_reduce_vc96;
      multm_reduce_sd98 <= multm_reduce_vc97;
      multm_reduce_sd99 <= multm_reduce_vc98;
      multm_reduce_sd100 <= multm_reduce_vc99;
      multm_reduce_sd101 <= multm_reduce_vc100;
      multm_reduce_sd102 <= multm_reduce_vc101;
      multm_reduce_sd103 <= multm_reduce_vc102;
      multm_reduce_sd104 <= multm_reduce_vc103;
      multm_reduce_sd105 <= multm_reduce_vc104;
      multm_reduce_sd106 <= multm_reduce_vc105;
      multm_reduce_sd107 <= multm_reduce_vc106;
      multm_reduce_sd108 <= multm_reduce_vc107;
      multm_reduce_sd109 <= multm_reduce_vc108;
      multm_reduce_sd110 <= multm_reduce_vc109;
      multm_reduce_sd111 <= multm_reduce_vc110;
      multm_reduce_sd112 <= multm_reduce_vc111;
      multm_reduce_sd113 <= multm_reduce_vc112;
      multm_reduce_sd114 <= multm_reduce_vc113;
      multm_reduce_sd115 <= multm_reduce_vc114;
      multm_reduce_sd116 <= multm_reduce_vc115;
      multm_reduce_sd117 <= multm_reduce_vc116;
      multm_reduce_sd118 <= multm_reduce_vc117;
      multm_reduce_sd119 <= multm_reduce_vc118;
      multm_reduce_sd120 <= multm_reduce_vc119;
      multm_reduce_sd121 <= multm_reduce_vc120;
      multm_reduce_sd122 <= multm_reduce_vc121;
      multm_reduce_sd123 <= multm_reduce_vc122;
      multm_reduce_sd124 <= multm_reduce_vc123;
      multm_reduce_sd125 <= multm_reduce_vc124;
      multm_reduce_sd126 <= multm_reduce_vc125;
      multm_reduce_sd127 <= multm_reduce_vc126;
      multm_reduce_sd128 <= multm_reduce_vc127;
      multm_reduce_sd129 <= multm_reduce_vc128;
      multm_reduce_sd130 <= multm_reduce_vc129;
      multm_reduce_sd131 <= multm_reduce_vc130;
      multm_reduce_sd132 <= multm_reduce_vc131;
      multm_reduce_sd133 <= multm_reduce_vc132;
      multm_reduce_sd134 <= multm_reduce_vc133;
      multm_reduce_sd135 <= multm_reduce_vc134;
      multm_reduce_sd136 <= multm_reduce_vc135;
      multm_reduce_sd137 <= multm_reduce_vc136;
      multm_reduce_sd138 <= multm_reduce_vc137;
      multm_reduce_sd139 <= multm_reduce_vc138;
      multm_reduce_sd140 <= multm_reduce_vc139;
      multm_reduce_sd141 <= multm_reduce_vc140;
      multm_reduce_sd142 <= multm_reduce_vc141;
      multm_reduce_sd143 <= multm_reduce_vc142;
      multm_reduce_sd144 <= multm_reduce_vc143;
      multm_reduce_sd145 <= multm_reduce_vc144;
      multm_reduce_sd146 <= multm_reduce_vc145;
      multm_reduce_sd147 <= multm_reduce_vc146;
      multm_reduce_sd148 <= multm_reduce_vc147;
      multm_reduce_sd149 <= multm_reduce_vc148;
      multm_reduce_sd150 <= multm_reduce_vc149;
      multm_reduce_sd151 <= multm_reduce_vc150;
      multm_reduce_sd152 <= multm_reduce_vc151;
      multm_reduce_sd153 <= multm_reduce_vc152;
      multm_reduce_sd154 <= multm_reduce_vc153;
      multm_reduce_sd155 <= multm_reduce_vc154;
      multm_reduce_sd156 <= multm_reduce_vc155;
      multm_reduce_sd157 <= multm_reduce_vc156;
      multm_reduce_sd158 <= multm_reduce_vc157;
      multm_reduce_sd159 <= multm_reduce_vc158;
      multm_reduce_sd160 <= multm_reduce_vc159;
      multm_reduce_sd161 <= multm_reduce_vc160;
      multm_reduce_sd162 <= multm_reduce_vc161;
      multm_reduce_sd163 <= multm_reduce_vc162;
      multm_reduce_sd164 <= multm_reduce_vc163;
      multm_reduce_sd165 <= multm_reduce_vc164;
      multm_reduce_sd166 <= multm_reduce_vc165;
      multm_reduce_sd167 <= multm_reduce_vc166;
      multm_reduce_sd168 <= multm_reduce_vc167;
      multm_reduce_sd169 <= multm_reduce_vc168;
      multm_reduce_sd170 <= multm_reduce_vc169;
      multm_reduce_sd171 <= multm_reduce_vc170;
      multm_reduce_sd172 <= multm_reduce_vc171;
      multm_reduce_sd173 <= multm_reduce_vc172;
      multm_reduce_sd174 <= multm_reduce_vc173;
      multm_reduce_sd175 <= multm_reduce_vc174;
      multm_reduce_sd176 <= multm_reduce_vc175;
      multm_reduce_sd177 <= multm_reduce_vc176;
      multm_reduce_sd178 <= multm_reduce_vc177;
      multm_reduce_sd179 <= multm_reduce_vc178;
      multm_reduce_sd180 <= multm_reduce_vc179;
      multm_reduce_sd181 <= multm_reduce_vc180;
      multm_reduce_sd182 <= multm_reduce_vc181;
      multm_reduce_sd183 <= multm_reduce_vc182;
      pipe0_x1 <= sa;
      pipe0_x2 <= pipe0_x1;
      pipe0_x3 <= pipe0_x2;
      pipe0_x4 <= pipe0_x3;
      pipe0_x5 <= pipe0_x4;
      pipe0_x6 <= pipe0_x5;
      pipe0_x7 <= pipe0_x6;
      pipe0_x8 <= pipe0_x7;
      pipe0_x9 <= pipe0_x8;
      pipe1_x1 <= sb;
      pipe1_x2 <= pipe1_x1;
      pipe1_x3 <= pipe1_x2;
      pipe1_x4 <= pipe1_x3;
      pipe1_x5 <= pipe1_x4;
      pipe1_x6 <= pipe1_x5;
      pipe1_x7 <= pipe1_x6;
      pipe1_x8 <= pipe1_x7;
      pipe1_x9 <= pipe1_x8;
      sa <= sar;
      sad <= pipe0_x9;
      sadd <= sad;
      sb <= sbr;
      sbd <= pipe1_x9;
      sbdd <= sbd;
      yc0_o <= pcr0;
      yc1_o <= pcr1;
      yc2_o <= pcr2;
      yc3_o <= pcr3;
      yc4_o <= pcr4;
      yc5_o <= pcr5;
      yc6_o <= pcr6;
      yc7_o <= pcr7;
      yc8_o <= pcr8;
      yc9_o <= pcr9;
      yc10_o <= pcr10;
      yc11_o <= pcr11;
      yc12_o <= pcr12;
      yc13_o <= pcr13;
      yc14_o <= pcr14;
      yc15_o <= pcr15;
      yc16_o <= pcr16;
      yc17_o <= pcr17;
      yc18_o <= pcr18;
      yc19_o <= pcr19;
      yc20_o <= pcr20;
      yc21_o <= pcr21;
      yc22_o <= pcr22;
      yc23_o <= pcr23;
      yc24_o <= pcr24;
      yc25_o <= pcr25;
      yc26_o <= pcr26;
      yc27_o <= pcr27;
      yc28_o <= pcr28;
      yc29_o <= pcr29;
      yc30_o <= pcr30;
      yc31_o <= pcr31;
      yc32_o <= pcr32;
      yc33_o <= pcr33;
      yc34_o <= pcr34;
      yc35_o <= pcr35;
      yc36_o <= pcr36;
      yc37_o <= pcr37;
      yc38_o <= pcr38;
      yc39_o <= pcr39;
      yc40_o <= pcr40;
      yc41_o <= pcr41;
      yc42_o <= pcr42;
      yc43_o <= pcr43;
      yc44_o <= pcr44;
      yc45_o <= pcr45;
      yc46_o <= pcr46;
      yc47_o <= pcr47;
      yc48_o <= pcr48;
      yc49_o <= pcr49;
      yc50_o <= pcr50;
      yc51_o <= pcr51;
      yc52_o <= pcr52;
      yc53_o <= pcr53;
      yc54_o <= pcr54;
      yc55_o <= pcr55;
      yc56_o <= pcr56;
      yc57_o <= pcr57;
      yc58_o <= pcr58;
      yc59_o <= pcr59;
      yc60_o <= pcr60;
      yc61_o <= pcr61;
      yc62_o <= pcr62;
      yc63_o <= pcr63;
      yc64_o <= pcr64;
      yc65_o <= pcr65;
      yc66_o <= pcr66;
      yc67_o <= pcr67;
      yc68_o <= pcr68;
      yc69_o <= pcr69;
      yc70_o <= pcr70;
      yc71_o <= pcr71;
      yc72_o <= pcr72;
      yc73_o <= pcr73;
      yc74_o <= pcr74;
      yc75_o <= pcr75;
      yc76_o <= pcr76;
      yc77_o <= pcr77;
      yc78_o <= pcr78;
      yc79_o <= pcr79;
      yc80_o <= pcr80;
      yc81_o <= pcr81;
      yc82_o <= pcr82;
      yc83_o <= pcr83;
      yc84_o <= pcr84;
      yc85_o <= pcr85;
      yc86_o <= pcr86;
      yc87_o <= pcr87;
      yc88_o <= pcr88;
      yc89_o <= pcr89;
      yc90_o <= pcr90;
      yc91_o <= pcr91;
      yc92_o <= pcr92;
      yc93_o <= pcr93;
      yc94_o <= pcr94;
      yc95_o <= pcr95;
      yc96_o <= pcr96;
      yc97_o <= pcr97;
      yc98_o <= pcr98;
      yc99_o <= pcr99;
      yc100_o <= pcr100;
      yc101_o <= pcr101;
      yc102_o <= pcr102;
      yc103_o <= pcr103;
      yc104_o <= pcr104;
      yc105_o <= pcr105;
      yc106_o <= pcr106;
      yc107_o <= pcr107;
      yc108_o <= pcr108;
      yc109_o <= pcr109;
      yc110_o <= pcr110;
      yc111_o <= pcr111;
      yc112_o <= pcr112;
      yc113_o <= pcr113;
      yc114_o <= pcr114;
      yc115_o <= pcr115;
      yc116_o <= pcr116;
      yc117_o <= pcr117;
      yc118_o <= pcr118;
      yc119_o <= pcr119;
      yc120_o <= pcr120;
      yc121_o <= pcr121;
      yc122_o <= pcr122;
      yc123_o <= pcr123;
      yc124_o <= pcr124;
      yc125_o <= pcr125;
      yc126_o <= pcr126;
      yc127_o <= pcr127;
      yc128_o <= pcr128;
      yc129_o <= pcr129;
      yc130_o <= pcr130;
      yc131_o <= pcr131;
      yc132_o <= pcr132;
      yc133_o <= pcr133;
      yc134_o <= pcr134;
      yc135_o <= pcr135;
      yc136_o <= pcr136;
      yc137_o <= pcr137;
      yc138_o <= pcr138;
      yc139_o <= pcr139;
      yc140_o <= pcr140;
      yc141_o <= pcr141;
      yc142_o <= pcr142;
      yc143_o <= pcr143;
      yc144_o <= pcr144;
      yc145_o <= pcr145;
      yc146_o <= pcr146;
      yc147_o <= pcr147;
      yc148_o <= pcr148;
      yc149_o <= pcr149;
      yc150_o <= pcr150;
      yc151_o <= pcr151;
      yc152_o <= pcr152;
      yc153_o <= pcr153;
      yc154_o <= pcr154;
      yc155_o <= pcr155;
      yc156_o <= pcr156;
      yc157_o <= pcr157;
      yc158_o <= pcr158;
      yc159_o <= pcr159;
      yc160_o <= pcr160;
      yc161_o <= pcr161;
      yc162_o <= pcr162;
      yc163_o <= pcr163;
      yc164_o <= pcr164;
      yc165_o <= pcr165;
      yc166_o <= pcr166;
      yc167_o <= pcr167;
      yc168_o <= pcr168;
      yc169_o <= pcr169;
      yc170_o <= pcr170;
      yc171_o <= pcr171;
      yc172_o <= pcr172;
      yc173_o <= pcr173;
      yc174_o <= pcr174;
      yc175_o <= pcr175;
      yc176_o <= pcr176;
      yc177_o <= pcr177;
      yc178_o <= pcr178;
      yc179_o <= pcr179;
      yc180_o <= pcr180;
      yc181_o <= pcr181;
      yc182_o <= pcr182;
      yc183_o <= pcr183;
      ys0_o <= psr0;
      ys1_o <= psr1;
      ys2_o <= psr2;
      ys3_o <= psr3;
      ys4_o <= psr4;
      ys5_o <= psr5;
      ys6_o <= psr6;
      ys7_o <= psr7;
      ys8_o <= psr8;
      ys9_o <= psr9;
      ys10_o <= psr10;
      ys11_o <= psr11;
      ys12_o <= psr12;
      ys13_o <= psr13;
      ys14_o <= psr14;
      ys15_o <= psr15;
      ys16_o <= psr16;
      ys17_o <= psr17;
      ys18_o <= psr18;
      ys19_o <= psr19;
      ys20_o <= psr20;
      ys21_o <= psr21;
      ys22_o <= psr22;
      ys23_o <= psr23;
      ys24_o <= psr24;
      ys25_o <= psr25;
      ys26_o <= psr26;
      ys27_o <= psr27;
      ys28_o <= psr28;
      ys29_o <= psr29;
      ys30_o <= psr30;
      ys31_o <= psr31;
      ys32_o <= psr32;
      ys33_o <= psr33;
      ys34_o <= psr34;
      ys35_o <= psr35;
      ys36_o <= psr36;
      ys37_o <= psr37;
      ys38_o <= psr38;
      ys39_o <= psr39;
      ys40_o <= psr40;
      ys41_o <= psr41;
      ys42_o <= psr42;
      ys43_o <= psr43;
      ys44_o <= psr44;
      ys45_o <= psr45;
      ys46_o <= psr46;
      ys47_o <= psr47;
      ys48_o <= psr48;
      ys49_o <= psr49;
      ys50_o <= psr50;
      ys51_o <= psr51;
      ys52_o <= psr52;
      ys53_o <= psr53;
      ys54_o <= psr54;
      ys55_o <= psr55;
      ys56_o <= psr56;
      ys57_o <= psr57;
      ys58_o <= psr58;
      ys59_o <= psr59;
      ys60_o <= psr60;
      ys61_o <= psr61;
      ys62_o <= psr62;
      ys63_o <= psr63;
      ys64_o <= psr64;
      ys65_o <= psr65;
      ys66_o <= psr66;
      ys67_o <= psr67;
      ys68_o <= psr68;
      ys69_o <= psr69;
      ys70_o <= psr70;
      ys71_o <= psr71;
      ys72_o <= psr72;
      ys73_o <= psr73;
      ys74_o <= psr74;
      ys75_o <= psr75;
      ys76_o <= psr76;
      ys77_o <= psr77;
      ys78_o <= psr78;
      ys79_o <= psr79;
      ys80_o <= psr80;
      ys81_o <= psr81;
      ys82_o <= psr82;
      ys83_o <= psr83;
      ys84_o <= psr84;
      ys85_o <= psr85;
      ys86_o <= psr86;
      ys87_o <= psr87;
      ys88_o <= psr88;
      ys89_o <= psr89;
      ys90_o <= psr90;
      ys91_o <= psr91;
      ys92_o <= psr92;
      ys93_o <= psr93;
      ys94_o <= psr94;
      ys95_o <= psr95;
      ys96_o <= psr96;
      ys97_o <= psr97;
      ys98_o <= psr98;
      ys99_o <= psr99;
      ys100_o <= psr100;
      ys101_o <= psr101;
      ys102_o <= psr102;
      ys103_o <= psr103;
      ys104_o <= psr104;
      ys105_o <= psr105;
      ys106_o <= psr106;
      ys107_o <= psr107;
      ys108_o <= psr108;
      ys109_o <= psr109;
      ys110_o <= psr110;
      ys111_o <= psr111;
      ys112_o <= psr112;
      ys113_o <= psr113;
      ys114_o <= psr114;
      ys115_o <= psr115;
      ys116_o <= psr116;
      ys117_o <= psr117;
      ys118_o <= psr118;
      ys119_o <= psr119;
      ys120_o <= psr120;
      ys121_o <= psr121;
      ys122_o <= psr122;
      ys123_o <= psr123;
      ys124_o <= psr124;
      ys125_o <= psr125;
      ys126_o <= psr126;
      ys127_o <= psr127;
      ys128_o <= psr128;
      ys129_o <= psr129;
      ys130_o <= psr130;
      ys131_o <= psr131;
      ys132_o <= psr132;
      ys133_o <= psr133;
      ys134_o <= psr134;
      ys135_o <= psr135;
      ys136_o <= psr136;
      ys137_o <= psr137;
      ys138_o <= psr138;
      ys139_o <= psr139;
      ys140_o <= psr140;
      ys141_o <= psr141;
      ys142_o <= psr142;
      ys143_o <= psr143;
      ys144_o <= psr144;
      ys145_o <= psr145;
      ys146_o <= psr146;
      ys147_o <= psr147;
      ys148_o <= psr148;
      ys149_o <= psr149;
      ys150_o <= psr150;
      ys151_o <= psr151;
      ys152_o <= psr152;
      ys153_o <= psr153;
      ys154_o <= psr154;
      ys155_o <= psr155;
      ys156_o <= psr156;
      ys157_o <= psr157;
      ys158_o <= psr158;
      ys159_o <= psr159;
      ys160_o <= psr160;
      ys161_o <= psr161;
      ys162_o <= psr162;
      ys163_o <= psr163;
      ys164_o <= psr164;
      ys165_o <= psr165;
      ys166_o <= psr166;
      ys167_o <= psr167;
      ys168_o <= psr168;
      ys169_o <= psr169;
      ys170_o <= psr170;
      ys171_o <= psr171;
      ys172_o <= psr172;
      ys173_o <= psr173;
      ys174_o <= psr174;
      ys175_o <= psr175;
      ys176_o <= psr176;
      ys177_o <= psr177;
      ys178_o <= psr178;
      ys179_o <= psr179;
      ys180_o <= psr180;
      ys181_o <= psr181;
      ys182_o <= psr182;
      ys183_o <= psr183;
    end

endmodule  // test_timelock_3

/*----------------------------------------------------------------------------+
| Primary inputs: 369                                                         |
| Primary outputs: 369                                                        |
| Registers: 2,321                                                            |
| Gates: 12,032                                                               |
| Fan-in: 25%=4 50%=6 75%=9 90%=9 95%=9 99%=9 max=9 (multm_qcp167)            |
| Fan-in cone: 25%=2 50%=9 75%=13 90%=17 95%=20 99%=20                        |
|   max=20 (multm_reduce_mulsc_mulb_cp181)                                    |
| Fan-out: 25%=2 50%=4 75%=7 90%=8 95%=8 99%=8 max=409 (sadd)                 |
| Duplication: 25%=1 50%=1 75%=1 90%=1 95%=1 99%=3 max=81 (sad)               |
| Fan-out load: 25%=2 50%=4 75%=7 90%=8 95%=8 99%=8                           |
|   max=8 (multm_reduce_sc25)                                                 |
+----------------------------------------------------------------------------*/
